module data_selector (clk, rst, wBusy, wSelec, wData, wRegs0, wRegs1, wRegs2, wRegs3, wRegs4, wRegs5, wRegs6, wRegs7, data_out);

input clk;
input rst;
input wBusy;
input [175:0] wSelec;
input [63:0] wData;
input [31:0] wRegs0;
input [31:0] wRegs1;
input [31:0] wRegs2;
input [31:0] wRegs3;
input [31:0] wRegs4;
input [31:0] wRegs5;
input [31:0] wRegs6;
input [31:0] wRegs7;
output [15:0] data_out;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX2 BUFX2_1 ( .A(clk), .Y(clk_hier0_bF_buf5) );
	BUFX2 BUFX2_2 ( .A(clk), .Y(clk_hier0_bF_buf4) );
	BUFX2 BUFX2_3 ( .A(clk), .Y(clk_hier0_bF_buf3) );
	BUFX2 BUFX2_4 ( .A(clk), .Y(clk_hier0_bF_buf2) );
	BUFX2 BUFX2_5 ( .A(clk), .Y(clk_hier0_bF_buf1) );
	BUFX2 BUFX2_6 ( .A(clk), .Y(clk_hier0_bF_buf0) );
	BUFX2 BUFX2_7 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf5) );
	BUFX2 BUFX2_8 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf4) );
	BUFX2 BUFX2_9 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf3) );
	BUFX2 BUFX2_10 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf2) );
	BUFX2 BUFX2_11 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf1) );
	BUFX2 BUFX2_12 ( .A(scheduler_block_scheduler_ctr_1_), .Y(scheduler_block_scheduler_ctr_1_bF_buf0) );
	BUFX4 BUFX4_1 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf42) );
	BUFX4 BUFX4_2 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf41) );
	BUFX4 BUFX4_3 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf40) );
	BUFX4 BUFX4_4 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf39) );
	BUFX4 BUFX4_5 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf38) );
	BUFX4 BUFX4_6 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf37) );
	BUFX4 BUFX4_7 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf36) );
	BUFX4 BUFX4_8 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf35) );
	BUFX4 BUFX4_9 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf34) );
	BUFX4 BUFX4_10 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf33) );
	BUFX4 BUFX4_11 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf32) );
	BUFX4 BUFX4_12 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf31) );
	BUFX4 BUFX4_13 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf30) );
	BUFX4 BUFX4_14 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf29) );
	BUFX4 BUFX4_15 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf28) );
	BUFX4 BUFX4_16 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf27) );
	BUFX4 BUFX4_17 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf26) );
	BUFX4 BUFX4_18 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf25) );
	BUFX4 BUFX4_19 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf24) );
	BUFX4 BUFX4_20 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf23) );
	BUFX4 BUFX4_21 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf22) );
	BUFX4 BUFX4_22 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf21) );
	BUFX4 BUFX4_23 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf20) );
	BUFX4 BUFX4_24 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf19) );
	BUFX4 BUFX4_25 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf18) );
	BUFX4 BUFX4_26 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf17) );
	BUFX4 BUFX4_27 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16) );
	BUFX4 BUFX4_28 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf15) );
	BUFX4 BUFX4_29 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf14) );
	BUFX4 BUFX4_30 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf13) );
	BUFX4 BUFX4_31 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf12) );
	BUFX4 BUFX4_32 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_33 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_34 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_35 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_36 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_37 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_38 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_39 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_40 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_41 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_42 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_43 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf0) );
	BUFX2 BUFX2_13 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf5) );
	BUFX2 BUFX2_14 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf4) );
	BUFX2 BUFX2_15 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf3) );
	BUFX2 BUFX2_16 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf2) );
	BUFX2 BUFX2_17 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf1) );
	BUFX2 BUFX2_18 ( .A(scheduler_block_scheduler_ctr_0_), .Y(scheduler_block_scheduler_ctr_0_bF_buf0) );
	BUFX2 BUFX2_19 ( .A(_8701_), .Y(_8701__bF_buf3) );
	BUFX2 BUFX2_20 ( .A(_8701_), .Y(_8701__bF_buf2) );
	BUFX2 BUFX2_21 ( .A(_8701_), .Y(_8701__bF_buf1) );
	BUFX2 BUFX2_22 ( .A(_8701_), .Y(_8701__bF_buf0) );
	BUFX2 BUFX2_23 ( .A(wBusy), .Y(wBusy_bF_buf4) );
	BUFX2 BUFX2_24 ( .A(wBusy), .Y(wBusy_bF_buf3) );
	BUFX2 BUFX2_25 ( .A(wBusy), .Y(wBusy_bF_buf2) );
	BUFX2 BUFX2_26 ( .A(wBusy), .Y(wBusy_bF_buf1) );
	BUFX2 BUFX2_27 ( .A(wBusy), .Y(wBusy_bF_buf0) );
	BUFX2 BUFX2_28 ( .A(rst), .Y(rst_bF_buf3) );
	BUFX2 BUFX2_29 ( .A(rst), .Y(rst_bF_buf2) );
	BUFX2 BUFX2_30 ( .A(rst), .Y(rst_bF_buf1) );
	BUFX2 BUFX2_31 ( .A(rst), .Y(rst_bF_buf0) );
	NAND2X1 NAND2X1_1 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_701_), .Y(_994_) );
	NAND2X1 NAND2X1_2 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_674_), .Y(_995_) );
	NAND2X1 NAND2X1_3 ( .A(_994_), .B(_995_), .Y(_996_) );
	INVX1 INVX1_1 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_997_) );
	NAND2X1 NAND2X1_4 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_673_), .Y(_998_) );
	OAI21X1 OAI21X1_1 ( .A(_997_), .B(_626_), .C(_998_), .Y(_999_) );
	NOR2X1 NOR2X1_1 ( .A(_996_), .B(_999_), .Y(_1000_) );
	NAND3X1 NAND3X1_1 ( .A(_990_), .B(_993_), .C(_1000_), .Y(_1001_) );
	NOR3X1 NOR3X1_1 ( .A(_988_), .B(_978_), .C(_1001_), .Y(_1002_) );
	INVX1 INVX1_2 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_1003_) );
	NAND2X1 NAND2X1_5 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_589_), .Y(_1004_) );
	OAI21X1 OAI21X1_2 ( .A(_594_), .B(_1003_), .C(_1004_), .Y(_1005_) );
	AOI21X1 AOI21X1_1 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_569_), .C(_1005_), .Y(_1006_) );
	INVX1 INVX1_3 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_1007_) );
	INVX1 INVX1_4 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_1008_) );
	OAI22X1 OAI22X1_1 ( .A(_913_), .B(_1008_), .C(_1007_), .D(_564_), .Y(_1009_) );
	INVX1 INVX1_5 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_1010_) );
	NAND2X1 NAND2X1_6 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_709_), .Y(_1011_) );
	OAI21X1 OAI21X1_3 ( .A(_574_), .B(_1010_), .C(_1011_), .Y(_1012_) );
	NOR2X1 NOR2X1_2 ( .A(_1012_), .B(_1009_), .Y(_1013_) );
	INVX1 INVX1_6 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_1014_) );
	INVX1 INVX1_7 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_1015_) );
	OAI22X1 OAI22X1_2 ( .A(_661_), .B(_1015_), .C(_1014_), .D(_662_), .Y(_1016_) );
	INVX1 INVX1_8 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_1017_) );
	NAND2X1 NAND2X1_7 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_708_), .Y(_1018_) );
	OAI21X1 OAI21X1_4 ( .A(_1017_), .B(_644_), .C(_1018_), .Y(_1019_) );
	NOR2X1 NOR2X1_3 ( .A(_1019_), .B(_1016_), .Y(_1020_) );
	NAND3X1 NAND3X1_2 ( .A(_1006_), .B(_1020_), .C(_1013_), .Y(_1021_) );
	AOI22X1 AOI22X1_1 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_666_), .C(_667_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_1022_) );
	AOI22X1 AOI22X1_2 ( .A(_669_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_670_), .Y(_1023_) );
	NAND2X1 NAND2X1_8 ( .A(_1022_), .B(_1023_), .Y(_1024_) );
	AOI22X1 AOI22X1_3 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_677_), .C(_676_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_1025_) );
	AOI22X1 AOI22X1_4 ( .A(_620_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_627_), .Y(_1026_) );
	NAND2X1 NAND2X1_9 ( .A(_1025_), .B(_1026_), .Y(_1027_) );
	NOR2X1 NOR2X1_4 ( .A(_1024_), .B(_1027_), .Y(_1028_) );
	AOI22X1 AOI22X1_5 ( .A(_681_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_682_), .Y(_1029_) );
	AOI22X1 AOI22X1_6 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_917_), .C(_684_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_1030_) );
	NAND2X1 NAND2X1_10 ( .A(_1030_), .B(_1029_), .Y(_1031_) );
	AOI22X1 AOI22X1_7 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_688_), .C(_689_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_1032_) );
	AOI22X1 AOI22X1_8 ( .A(_691_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_692_), .Y(_1033_) );
	NAND2X1 NAND2X1_11 ( .A(_1033_), .B(_1032_), .Y(_1034_) );
	NOR2X1 NOR2X1_5 ( .A(_1031_), .B(_1034_), .Y(_1035_) );
	NAND2X1 NAND2X1_12 ( .A(_1035_), .B(_1028_), .Y(_1036_) );
	AOI22X1 AOI22X1_9 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_698_), .C(_599_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_1037_) );
	AOI22X1 AOI22X1_10 ( .A(_622_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_700_), .Y(_1038_) );
	NAND2X1 NAND2X1_13 ( .A(_1037_), .B(_1038_), .Y(_1039_) );
	AOI22X1 AOI22X1_11 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_706_), .C(_704_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_1040_) );
	AOI22X1 AOI22X1_12 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_636_), .C(_685_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_1041_) );
	NAND2X1 NAND2X1_14 ( .A(_1041_), .B(_1040_), .Y(_1042_) );
	NOR2X1 NOR2X1_6 ( .A(_1042_), .B(_1039_), .Y(_1043_) );
	AOI22X1 AOI22X1_13 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_713_), .C(_714_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_1044_) );
	NAND2X1 NAND2X1_15 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_716_), .Y(_1045_) );
	NAND2X1 NAND2X1_16 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_718_), .Y(_1046_) );
	NAND3X1 NAND3X1_3 ( .A(_1045_), .B(_1046_), .C(_1044_), .Y(_1047_) );
	AOI22X1 AOI22X1_14 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_722_), .C(_721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_1048_) );
	AOI22X1 AOI22X1_15 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_725_), .C(_724_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_1049_) );
	NAND2X1 NAND2X1_17 ( .A(_1048_), .B(_1049_), .Y(_1050_) );
	NOR2X1 NOR2X1_7 ( .A(_1050_), .B(_1047_), .Y(_1051_) );
	NAND2X1 NAND2X1_18 ( .A(_1043_), .B(_1051_), .Y(_1052_) );
	NOR3X1 NOR3X1_2 ( .A(_1036_), .B(_1021_), .C(_1052_), .Y(_1053_) );
	NAND2X1 NAND2X1_19 ( .A(wData[59]), .B(_755_), .Y(_1054_) );
	OAI21X1 OAI21X1_5 ( .A(_539_), .B(wBusy_bF_buf4), .C(_1054_), .Y(_1055_) );
	NAND2X1 NAND2X1_20 ( .A(wData[7]), .B(_746_), .Y(_1056_) );
	NAND2X1 NAND2X1_21 ( .A(wData[55]), .B(_756_), .Y(_1057_) );
	AOI22X1 AOI22X1_16 ( .A(wData[63]), .B(_758_), .C(_748_), .D(wData[31]), .Y(_1058_) );
	NAND3X1 NAND3X1_4 ( .A(_1056_), .B(_1057_), .C(_1058_), .Y(_1059_) );
	OR2X2 OR2X2_1 ( .A(_1059_), .B(_1055_), .Y(_1060_) );
	INVX1 INVX1_9 ( .A(wData[51]), .Y(_1061_) );
	NAND2X1 NAND2X1_22 ( .A(wData[47]), .B(_759_), .Y(_1062_) );
	OAI21X1 OAI21X1_6 ( .A(_1061_), .B(_771_), .C(_1062_), .Y(_1063_) );
	AOI21X1 AOI21X1_2 ( .A(wData[3]), .B(_766_), .C(_1063_), .Y(_1064_) );
	AOI22X1 AOI22X1_17 ( .A(_772_), .B(wData[11]), .C(wData[15]), .D(_773_), .Y(_1065_) );
	AOI22X1 AOI22X1_18 ( .A(_735_), .B(wData[23]), .C(wData[27]), .D(_742_), .Y(_1066_) );
	AND2X2 AND2X2_1 ( .A(_1065_), .B(_1066_), .Y(_1067_) );
	NAND2X1 NAND2X1_23 ( .A(wData[39]), .B(_764_), .Y(_1068_) );
	NAND2X1 NAND2X1_24 ( .A(wData[43]), .B(_762_), .Y(_1069_) );
	NAND2X1 NAND2X1_25 ( .A(_1068_), .B(_1069_), .Y(_1070_) );
	NAND2X1 NAND2X1_26 ( .A(wData[19]), .B(_738_), .Y(_1071_) );
	NAND2X1 NAND2X1_27 ( .A(wData[35]), .B(_752_), .Y(_1072_) );
	NAND2X1 NAND2X1_28 ( .A(_1071_), .B(_1072_), .Y(_1073_) );
	NOR2X1 NOR2X1_8 ( .A(_1070_), .B(_1073_), .Y(_1074_) );
	NAND3X1 NAND3X1_5 ( .A(_1067_), .B(_1064_), .C(_1074_), .Y(_1075_) );
	NOR2X1 NOR2X1_9 ( .A(_1060_), .B(_1075_), .Y(_1076_) );
	AOI21X1 AOI21X1_3 ( .A(_1002_), .B(_1053_), .C(_1076_), .Y(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_3_) );
	INVX1 INVX1_10 ( .A(wSelec[22]), .Y(_1077_) );
	NOR2X1 NOR2X1_10 ( .A(wBusy_bF_buf3), .B(_1077_), .Y(_1078_) );
	INVX1 INVX1_11 ( .A(_1078_), .Y(_1079_) );
	INVX1 INVX1_12 ( .A(wSelec[32]), .Y(_1080_) );
	NAND2X1 NAND2X1_29 ( .A(wSelec[31]), .B(_1080_), .Y(_1081_) );
	INVX2 INVX2_1 ( .A(_1081_), .Y(_1082_) );
	OR2X2 OR2X2_2 ( .A(wSelec[28]), .B(wSelec[27]), .Y(_1083_) );
	INVX1 INVX1_13 ( .A(wSelec[30]), .Y(_1084_) );
	NAND2X1 NAND2X1_30 ( .A(wSelec[29]), .B(_1084_), .Y(_1085_) );
	NOR2X1 NOR2X1_11 ( .A(_1083_), .B(_1085_), .Y(_1086_) );
	AND2X2 AND2X2_2 ( .A(_1086_), .B(_1082_), .Y(_1087_) );
	AOI21X1 AOI21X1_4 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_1087_), .C(_1079_), .Y(_1088_) );
	INVX1 INVX1_14 ( .A(wSelec[28]), .Y(_1089_) );
	NAND2X1 NAND2X1_31 ( .A(wSelec[27]), .B(_1089_), .Y(_1090_) );
	OR2X2 OR2X2_3 ( .A(wSelec[29]), .B(wSelec[30]), .Y(_1091_) );
	NOR2X1 NOR2X1_12 ( .A(_1091_), .B(_1090_), .Y(_1092_) );
	NAND2X1 NAND2X1_32 ( .A(_1082_), .B(_1092_), .Y(_1093_) );
	INVX1 INVX1_15 ( .A(_1093_), .Y(_1094_) );
	INVX1 INVX1_16 ( .A(wSelec[27]), .Y(_1095_) );
	NAND2X1 NAND2X1_33 ( .A(wSelec[28]), .B(_1095_), .Y(_1096_) );
	INVX1 INVX1_17 ( .A(wSelec[29]), .Y(_1097_) );
	NAND2X1 NAND2X1_34 ( .A(wSelec[30]), .B(_1097_), .Y(_1098_) );
	NOR2X1 NOR2X1_13 ( .A(_1096_), .B(_1098_), .Y(_1099_) );
	NAND2X1 NAND2X1_35 ( .A(wSelec[31]), .B(wSelec[32]), .Y(_1100_) );
	INVX1 INVX1_18 ( .A(_1100_), .Y(_1101_) );
	NAND2X1 NAND2X1_36 ( .A(_1101_), .B(_1099_), .Y(_1102_) );
	INVX1 INVX1_19 ( .A(_1102_), .Y(_1103_) );
	AOI22X1 AOI22X1_19 ( .A(_1094_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_1103_), .Y(_1104_) );
	OR2X2 OR2X2_4 ( .A(_1090_), .B(_1091_), .Y(_1105_) );
	OR2X2 OR2X2_5 ( .A(wSelec[31]), .B(wSelec[32]), .Y(_1106_) );
	NOR2X1 NOR2X1_14 ( .A(_1106_), .B(_1105_), .Y(_1107_) );
	NOR2X1 NOR2X1_15 ( .A(_1085_), .B(_1090_), .Y(_1108_) );
	INVX1 INVX1_20 ( .A(wSelec[31]), .Y(_1109_) );
	NAND2X1 NAND2X1_37 ( .A(wSelec[32]), .B(_1109_), .Y(_1110_) );
	INVX2 INVX2_2 ( .A(_1110_), .Y(_1111_) );
	NAND2X1 NAND2X1_38 ( .A(_1111_), .B(_1108_), .Y(_1112_) );
	INVX1 INVX1_21 ( .A(_1112_), .Y(_1113_) );
	AOI22X1 AOI22X1_20 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_1107_), .C(_1113_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_1114_) );
	NAND3X1 NAND3X1_6 ( .A(_1088_), .B(_1114_), .C(_1104_), .Y(_1115_) );
	NOR2X1 NOR2X1_16 ( .A(wSelec[28]), .B(wSelec[27]), .Y(_1116_) );
	NOR2X1 NOR2X1_17 ( .A(wSelec[29]), .B(wSelec[30]), .Y(_1117_) );
	NAND2X1 NAND2X1_39 ( .A(_1116_), .B(_1117_), .Y(_1118_) );
	NOR2X1 NOR2X1_18 ( .A(_1081_), .B(_1118_), .Y(_1119_) );
	NAND2X1 NAND2X1_40 ( .A(wSelec[28]), .B(wSelec[27]), .Y(_1120_) );
	NOR3X1 NOR3X1_3 ( .A(_1091_), .B(_1120_), .C(_1081_), .Y(_1121_) );
	AOI22X1 AOI22X1_21 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_1121_), .C(_1119_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_1122_) );
	INVX1 INVX1_22 ( .A(_1106_), .Y(_1123_) );
	NOR2X1 NOR2X1_19 ( .A(_1091_), .B(_1096_), .Y(_1124_) );
	AND2X2 AND2X2_3 ( .A(_1124_), .B(_1123_), .Y(_1125_) );
	NAND2X1 NAND2X1_41 ( .A(wSelec[29]), .B(wSelec[30]), .Y(_1126_) );
	NOR3X1 NOR3X1_4 ( .A(_1100_), .B(_1120_), .C(_1126_), .Y(_1127_) );
	AOI22X1 AOI22X1_22 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_1127_), .C(_1125_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_1128_) );
	INVX1 INVX1_23 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_1129_) );
	INVX1 INVX1_24 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_1130_) );
	NOR2X1 NOR2X1_20 ( .A(_1090_), .B(_1098_), .Y(_1131_) );
	NAND2X1 NAND2X1_42 ( .A(_1101_), .B(_1131_), .Y(_1132_) );
	NOR2X1 NOR2X1_21 ( .A(_1120_), .B(_1126_), .Y(_1133_) );
	NAND2X1 NAND2X1_43 ( .A(_1133_), .B(_1111_), .Y(_1134_) );
	OAI22X1 OAI22X1_3 ( .A(_1129_), .B(_1134_), .C(_1132_), .D(_1130_), .Y(_1135_) );
	INVX1 INVX1_25 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_1136_) );
	NOR3X1 NOR3X1_5 ( .A(_1081_), .B(_1096_), .C(_1098_), .Y(_1137_) );
	NAND2X1 NAND2X1_44 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_1137_), .Y(_1138_) );
	NOR2X1 NOR2X1_22 ( .A(_1120_), .B(_1085_), .Y(_1139_) );
	NAND2X1 NAND2X1_45 ( .A(_1111_), .B(_1139_), .Y(_1140_) );
	OAI21X1 OAI21X1_7 ( .A(_1136_), .B(_1140_), .C(_1138_), .Y(_1141_) );
	NOR2X1 NOR2X1_23 ( .A(_1135_), .B(_1141_), .Y(_1142_) );
	NAND3X1 NAND3X1_7 ( .A(_1122_), .B(_1128_), .C(_1142_), .Y(_1143_) );
	INVX1 INVX1_26 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_1144_) );
	INVX1 INVX1_27 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_1145_) );
	NOR2X1 NOR2X1_24 ( .A(_1085_), .B(_1096_), .Y(_1146_) );
	NAND2X1 NAND2X1_46 ( .A(_1082_), .B(_1146_), .Y(_1147_) );
	NOR2X1 NOR2X1_25 ( .A(_1083_), .B(_1098_), .Y(_1148_) );
	NAND2X1 NAND2X1_47 ( .A(_1082_), .B(_1148_), .Y(_1149_) );
	OAI22X1 OAI22X1_4 ( .A(_1149_), .B(_1144_), .C(_1145_), .D(_1147_), .Y(_1150_) );
	INVX1 INVX1_28 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_1151_) );
	INVX1 INVX1_29 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_1152_) );
	NAND2X1 NAND2X1_48 ( .A(_1111_), .B(_1146_), .Y(_1153_) );
	NOR2X1 NOR2X1_26 ( .A(_1120_), .B(_1091_), .Y(_1154_) );
	NAND2X1 NAND2X1_49 ( .A(_1111_), .B(_1154_), .Y(_1155_) );
	OAI22X1 OAI22X1_5 ( .A(_1151_), .B(_1155_), .C(_1153_), .D(_1152_), .Y(_1156_) );
	NOR2X1 NOR2X1_27 ( .A(_1156_), .B(_1150_), .Y(_1157_) );
	NOR3X1 NOR3X1_6 ( .A(_1090_), .B(_1126_), .C(_1110_), .Y(_1158_) );
	NAND2X1 NAND2X1_50 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_1158_), .Y(_1159_) );
	NOR3X1 NOR3X1_7 ( .A(_1098_), .B(_1120_), .C(_1110_), .Y(_1160_) );
	NAND2X1 NAND2X1_51 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_1160_), .Y(_1161_) );
	NAND2X1 NAND2X1_52 ( .A(_1159_), .B(_1161_), .Y(_1162_) );
	INVX1 INVX1_30 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_1163_) );
	NAND2X1 NAND2X1_53 ( .A(_1101_), .B(_1086_), .Y(_1164_) );
	NOR3X1 NOR3X1_8 ( .A(_1096_), .B(_1098_), .C(_1110_), .Y(_1165_) );
	NAND2X1 NAND2X1_54 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_1165_), .Y(_1166_) );
	OAI21X1 OAI21X1_8 ( .A(_1163_), .B(_1164_), .C(_1166_), .Y(_1167_) );
	NOR2X1 NOR2X1_28 ( .A(_1162_), .B(_1167_), .Y(_1168_) );
	NAND2X1 NAND2X1_55 ( .A(_1157_), .B(_1168_), .Y(_1169_) );
	NOR3X1 NOR3X1_9 ( .A(_1115_), .B(_1169_), .C(_1143_), .Y(_1170_) );
	NAND2X1 NAND2X1_56 ( .A(_1082_), .B(_1139_), .Y(_1171_) );
	INVX1 INVX1_31 ( .A(_1171_), .Y(_1172_) );
	INVX1 INVX1_32 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_1173_) );
	NOR3X1 NOR3X1_10 ( .A(_1083_), .B(_1106_), .C(_1085_), .Y(_1174_) );
	NAND2X1 NAND2X1_57 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_1174_), .Y(_1175_) );
	NAND2X1 NAND2X1_58 ( .A(_1123_), .B(_1146_), .Y(_1176_) );
	OAI21X1 OAI21X1_9 ( .A(_1176_), .B(_1173_), .C(_1175_), .Y(_1177_) );
	AOI21X1 AOI21X1_5 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_1172_), .C(_1177_), .Y(_1178_) );
	INVX1 INVX1_33 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_1179_) );
	INVX1 INVX1_34 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_1180_) );
	NOR2X1 NOR2X1_29 ( .A(_1126_), .B(_1083_), .Y(_1181_) );
	NAND2X1 NAND2X1_59 ( .A(_1082_), .B(_1181_), .Y(_1182_) );
	NAND2X1 NAND2X1_60 ( .A(_1123_), .B(_1108_), .Y(_1183_) );
	OAI22X1 OAI22X1_6 ( .A(_1180_), .B(_1182_), .C(_1183_), .D(_1179_), .Y(_1184_) );
	INVX1 INVX1_35 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_1185_) );
	INVX1 INVX1_36 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_1186_) );
	NAND2X1 NAND2X1_61 ( .A(_1082_), .B(_1108_), .Y(_1187_) );
	NAND2X1 NAND2X1_62 ( .A(_1123_), .B(_1154_), .Y(_1188_) );
	OAI22X1 OAI22X1_7 ( .A(_1185_), .B(_1188_), .C(_1187_), .D(_1186_), .Y(_1189_) );
	NOR2X1 NOR2X1_30 ( .A(_1184_), .B(_1189_), .Y(_1190_) );
	INVX1 INVX1_37 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_1191_) );
	NOR3X1 NOR3X1_11 ( .A(_1106_), .B(_1120_), .C(_1085_), .Y(_1192_) );
	NAND2X1 NAND2X1_63 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_1192_), .Y(_1193_) );
	OR2X2 OR2X2_6 ( .A(_1118_), .B(_1100_), .Y(_1194_) );
	OAI21X1 OAI21X1_10 ( .A(_1191_), .B(_1194_), .C(_1193_), .Y(_1195_) );
	INVX1 INVX1_38 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_1196_) );
	INVX1 INVX1_39 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_1197_) );
	NOR2X1 NOR2X1_31 ( .A(_1126_), .B(_1096_), .Y(_1198_) );
	NAND2X1 NAND2X1_64 ( .A(_1082_), .B(_1198_), .Y(_1199_) );
	NAND2X1 NAND2X1_65 ( .A(_1101_), .B(_1092_), .Y(_1200_) );
	OAI22X1 OAI22X1_8 ( .A(_1199_), .B(_1197_), .C(_1196_), .D(_1200_), .Y(_1201_) );
	NOR2X1 NOR2X1_32 ( .A(_1195_), .B(_1201_), .Y(_1202_) );
	NAND3X1 NAND3X1_8 ( .A(_1178_), .B(_1202_), .C(_1190_), .Y(_1203_) );
	NOR3X1 NOR3X1_12 ( .A(_1083_), .B(_1091_), .C(_1106_), .Y(_1204_) );
	NOR3X1 NOR3X1_13 ( .A(_1100_), .B(_1126_), .C(_1090_), .Y(_1205_) );
	AOI22X1 AOI22X1_23 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_1204_), .C(_1205_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_1206_) );
	NOR3X1 NOR3X1_14 ( .A(_1100_), .B(_1126_), .C(_1096_), .Y(_1207_) );
	NOR3X1 NOR3X1_15 ( .A(_1100_), .B(_1120_), .C(_1098_), .Y(_1208_) );
	AOI22X1 AOI22X1_24 ( .A(_1207_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_1208_), .Y(_1209_) );
	NAND2X1 NAND2X1_66 ( .A(_1206_), .B(_1209_), .Y(_1210_) );
	NOR3X1 NOR3X1_16 ( .A(_1098_), .B(_1083_), .C(_1110_), .Y(_1211_) );
	NOR3X1 NOR3X1_17 ( .A(_1090_), .B(_1098_), .C(_1110_), .Y(_1212_) );
	AOI22X1 AOI22X1_25 ( .A(_1211_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_1212_), .Y(_1213_) );
	NOR3X1 NOR3X1_18 ( .A(_1081_), .B(_1126_), .C(_1090_), .Y(_1214_) );
	NOR3X1 NOR3X1_19 ( .A(_1120_), .B(_1126_), .C(_1081_), .Y(_1215_) );
	AOI22X1 AOI22X1_26 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_1215_), .C(_1214_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_1216_) );
	NAND2X1 NAND2X1_67 ( .A(_1216_), .B(_1213_), .Y(_1217_) );
	NOR2X1 NOR2X1_33 ( .A(_1210_), .B(_1217_), .Y(_1218_) );
	NOR3X1 NOR3X1_20 ( .A(_1106_), .B(_1126_), .C(_1090_), .Y(_1219_) );
	NOR3X1 NOR3X1_21 ( .A(_1106_), .B(_1126_), .C(_1096_), .Y(_1220_) );
	AOI22X1 AOI22X1_27 ( .A(_1219_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_1220_), .Y(_1221_) );
	NOR3X1 NOR3X1_22 ( .A(_1106_), .B(_1120_), .C(_1098_), .Y(_1222_) );
	NOR3X1 NOR3X1_23 ( .A(_1081_), .B(_1091_), .C(_1096_), .Y(_1223_) );
	AOI22X1 AOI22X1_28 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_1222_), .C(_1223_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_1224_) );
	NAND2X1 NAND2X1_68 ( .A(_1221_), .B(_1224_), .Y(_1225_) );
	NOR3X1 NOR3X1_24 ( .A(_1120_), .B(_1126_), .C(_1106_), .Y(_1226_) );
	NOR3X1 NOR3X1_25 ( .A(_1096_), .B(_1091_), .C(_1110_), .Y(_1227_) );
	AOI22X1 AOI22X1_29 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_1226_), .C(_1227_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_1228_) );
	NOR3X1 NOR3X1_26 ( .A(_1083_), .B(_1091_), .C(_1110_), .Y(_1229_) );
	NOR3X1 NOR3X1_27 ( .A(_1083_), .B(_1126_), .C(_1110_), .Y(_1230_) );
	AOI22X1 AOI22X1_30 ( .A(_1229_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_1230_), .Y(_1231_) );
	NAND2X1 NAND2X1_69 ( .A(_1231_), .B(_1228_), .Y(_1232_) );
	NOR2X1 NOR2X1_34 ( .A(_1225_), .B(_1232_), .Y(_1233_) );
	NAND2X1 NAND2X1_70 ( .A(_1233_), .B(_1218_), .Y(_1234_) );
	NOR3X1 NOR3X1_28 ( .A(_1081_), .B(_1120_), .C(_1098_), .Y(_1235_) );
	NOR3X1 NOR3X1_29 ( .A(_1091_), .B(_1100_), .C(_1096_), .Y(_1236_) );
	AOI22X1 AOI22X1_31 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_1236_), .C(_1235_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_1237_) );
	NOR3X1 NOR3X1_30 ( .A(_1085_), .B(_1083_), .C(_1110_), .Y(_1238_) );
	NOR3X1 NOR3X1_31 ( .A(_1096_), .B(_1126_), .C(_1110_), .Y(_1239_) );
	AOI22X1 AOI22X1_32 ( .A(_1238_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_1239_), .Y(_1240_) );
	NAND2X1 NAND2X1_71 ( .A(_1237_), .B(_1240_), .Y(_1241_) );
	NOR3X1 NOR3X1_32 ( .A(_1081_), .B(_1090_), .C(_1098_), .Y(_1242_) );
	NAND2X1 NAND2X1_72 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_1242_), .Y(_1243_) );
	NOR3X1 NOR3X1_33 ( .A(_1100_), .B(_1120_), .C(_1085_), .Y(_1244_) );
	NAND2X1 NAND2X1_73 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_1244_), .Y(_1245_) );
	NOR3X1 NOR3X1_34 ( .A(_1083_), .B(_1126_), .C(_1106_), .Y(_1246_) );
	NOR3X1 NOR3X1_35 ( .A(_1083_), .B(_1100_), .C(_1098_), .Y(_1247_) );
	AOI22X1 AOI22X1_33 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_1246_), .C(_1247_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_1248_) );
	NAND3X1 NAND3X1_9 ( .A(_1243_), .B(_1245_), .C(_1248_), .Y(_1249_) );
	NOR2X1 NOR2X1_35 ( .A(_1249_), .B(_1241_), .Y(_1250_) );
	NOR3X1 NOR3X1_36 ( .A(_1083_), .B(_1106_), .C(_1098_), .Y(_1251_) );
	NOR3X1 NOR3X1_37 ( .A(_1085_), .B(_1100_), .C(_1090_), .Y(_1252_) );
	AOI22X1 AOI22X1_34 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_1251_), .C(_1252_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_1253_) );
	NOR3X1 NOR3X1_38 ( .A(_1085_), .B(_1100_), .C(_1096_), .Y(_1254_) );
	NAND2X1 NAND2X1_74 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_1254_), .Y(_1255_) );
	NOR3X1 NOR3X1_39 ( .A(_1090_), .B(_1091_), .C(_1110_), .Y(_1256_) );
	NAND2X1 NAND2X1_75 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_1256_), .Y(_1257_) );
	NAND3X1 NAND3X1_10 ( .A(_1255_), .B(_1257_), .C(_1253_), .Y(_1258_) );
	NOR3X1 NOR3X1_40 ( .A(_1090_), .B(_1106_), .C(_1098_), .Y(_1259_) );
	NOR3X1 NOR3X1_41 ( .A(_1100_), .B(_1126_), .C(_1083_), .Y(_1260_) );
	AOI22X1 AOI22X1_35 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_1260_), .C(_1259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_1261_) );
	NOR3X1 NOR3X1_42 ( .A(_1096_), .B(_1106_), .C(_1098_), .Y(_1262_) );
	NOR3X1 NOR3X1_43 ( .A(_1100_), .B(_1120_), .C(_1091_), .Y(_1263_) );
	AOI22X1 AOI22X1_36 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_1263_), .C(_1262_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_1264_) );
	NAND2X1 NAND2X1_76 ( .A(_1261_), .B(_1264_), .Y(_1265_) );
	NOR2X1 NOR2X1_36 ( .A(_1265_), .B(_1258_), .Y(_1266_) );
	NAND2X1 NAND2X1_77 ( .A(_1250_), .B(_1266_), .Y(_1267_) );
	NOR3X1 NOR3X1_44 ( .A(_1234_), .B(_1203_), .C(_1267_), .Y(_1268_) );
	INVX1 INVX1_40 ( .A(wSelec[24]), .Y(_1269_) );
	NAND2X1 NAND2X1_78 ( .A(wSelec[23]), .B(_1269_), .Y(_1270_) );
	INVX1 INVX1_41 ( .A(wSelec[26]), .Y(_1271_) );
	NAND2X1 NAND2X1_79 ( .A(wSelec[25]), .B(_1271_), .Y(_1272_) );
	NOR2X1 NOR2X1_37 ( .A(_1270_), .B(_1272_), .Y(_1273_) );
	NOR2X1 NOR2X1_38 ( .A(wSelec[24]), .B(wSelec[23]), .Y(_1274_) );
	INVX1 INVX1_42 ( .A(_1274_), .Y(_1275_) );
	NOR2X1 NOR2X1_39 ( .A(_1272_), .B(_1275_), .Y(_1276_) );
	AOI22X1 AOI22X1_37 ( .A(wData[20]), .B(_1273_), .C(_1276_), .D(wData[16]), .Y(_1277_) );
	INVX1 INVX1_43 ( .A(wSelec[23]), .Y(_1278_) );
	NAND2X1 NAND2X1_80 ( .A(wSelec[24]), .B(_1278_), .Y(_1279_) );
	NOR2X1 NOR2X1_40 ( .A(_1279_), .B(_1272_), .Y(_1280_) );
	NAND2X1 NAND2X1_81 ( .A(wData[24]), .B(_1280_), .Y(_1281_) );
	INVX1 INVX1_44 ( .A(wSelec[25]), .Y(_1282_) );
	NAND2X1 NAND2X1_82 ( .A(_1282_), .B(_1271_), .Y(_1283_) );
	NOR2X1 NOR2X1_41 ( .A(_1270_), .B(_1283_), .Y(_1284_) );
	NAND2X1 NAND2X1_83 ( .A(wSelec[24]), .B(wSelec[23]), .Y(_1285_) );
	NOR2X1 NOR2X1_42 ( .A(_1285_), .B(_1272_), .Y(_1286_) );
	AOI22X1 AOI22X1_38 ( .A(_1286_), .B(wData[28]), .C(wData[4]), .D(_1284_), .Y(_1287_) );
	NAND3X1 NAND3X1_11 ( .A(_1281_), .B(_1287_), .C(_1277_), .Y(_1288_) );
	NAND2X1 NAND2X1_84 ( .A(wSelec[26]), .B(_1282_), .Y(_1289_) );
	NOR2X1 NOR2X1_43 ( .A(_1289_), .B(_1275_), .Y(_1290_) );
	NAND2X1 NAND2X1_85 ( .A(wData[32]), .B(_1290_), .Y(_1291_) );
	NAND2X1 NAND2X1_86 ( .A(wSelec[25]), .B(wSelec[26]), .Y(_1292_) );
	NOR2X1 NOR2X1_44 ( .A(_1292_), .B(_1279_), .Y(_1293_) );
	NOR2X1 NOR2X1_45 ( .A(_1292_), .B(_1270_), .Y(_1294_) );
	AOI22X1 AOI22X1_39 ( .A(_1293_), .B(wData[56]), .C(wData[52]), .D(_1294_), .Y(_1295_) );
	NOR2X1 NOR2X1_46 ( .A(_1285_), .B(_1292_), .Y(_1296_) );
	NOR2X1 NOR2X1_47 ( .A(_1285_), .B(_1289_), .Y(_1297_) );
	AOI22X1 AOI22X1_40 ( .A(wData[60]), .B(_1296_), .C(_1297_), .D(wData[44]), .Y(_1298_) );
	NAND3X1 NAND3X1_12 ( .A(_1291_), .B(_1298_), .C(_1295_), .Y(_1299_) );
	NOR2X1 NOR2X1_48 ( .A(_1279_), .B(_1289_), .Y(_1300_) );
	NAND2X1 NAND2X1_87 ( .A(wData[40]), .B(_1300_), .Y(_1301_) );
	NOR2X1 NOR2X1_49 ( .A(_1289_), .B(_1270_), .Y(_1302_) );
	NAND2X1 NAND2X1_88 ( .A(wData[36]), .B(_1302_), .Y(_1303_) );
	NOR2X1 NOR2X1_50 ( .A(_1283_), .B(_1275_), .Y(_1304_) );
	NAND2X1 NAND2X1_89 ( .A(wData[0]), .B(_1304_), .Y(_1305_) );
	NAND3X1 NAND3X1_13 ( .A(_1301_), .B(_1303_), .C(_1305_), .Y(_1306_) );
	INVX1 INVX1_45 ( .A(wData[48]), .Y(_1307_) );
	NOR2X1 NOR2X1_51 ( .A(_1282_), .B(_1271_), .Y(_1308_) );
	NAND2X1 NAND2X1_90 ( .A(_1274_), .B(_1308_), .Y(_1309_) );
	NOR2X1 NOR2X1_52 ( .A(_1279_), .B(_1283_), .Y(_1310_) );
	NOR2X1 NOR2X1_53 ( .A(_1285_), .B(_1283_), .Y(_1311_) );
	AOI22X1 AOI22X1_41 ( .A(_1310_), .B(wData[8]), .C(wData[12]), .D(_1311_), .Y(_1312_) );
	OAI21X1 OAI21X1_11 ( .A(_1307_), .B(_1309_), .C(_1312_), .Y(_1313_) );
	OR2X2 OR2X2_7 ( .A(_1313_), .B(_1306_), .Y(_1314_) );
	NOR3X1 NOR3X1_45 ( .A(_1288_), .B(_1299_), .C(_1314_), .Y(_1315_) );
	AND2X2 AND2X2_4 ( .A(_1315_), .B(_1079_), .Y(_1316_) );
	AOI21X1 AOI21X1_6 ( .A(_1170_), .B(_1268_), .C(_1316_), .Y(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_0_) );
	INVX1 INVX1_46 ( .A(_1187_), .Y(_1317_) );
	AOI21X1 AOI21X1_7 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_1317_), .C(_1079_), .Y(_1318_) );
	AOI22X1 AOI22X1_42 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_1087_), .C(_1103_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_1319_) );
	AOI22X1 AOI22X1_43 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_1107_), .C(_1113_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_1320_) );
	NAND3X1 NAND3X1_14 ( .A(_1318_), .B(_1319_), .C(_1320_), .Y(_1321_) );
	INVX1 INVX1_47 ( .A(_1147_), .Y(_1322_) );
	AOI22X1 AOI22X1_44 ( .A(_1172_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_1322_), .Y(_1323_) );
	AOI22X1 AOI22X1_45 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_1246_), .C(_1125_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_1324_) );
	INVX1 INVX1_48 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_1325_) );
	INVX1 INVX1_49 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_1326_) );
	OAI22X1 OAI22X1_9 ( .A(_1325_), .B(_1134_), .C(_1132_), .D(_1326_), .Y(_1327_) );
	INVX1 INVX1_50 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_1328_) );
	NAND2X1 NAND2X1_91 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_1235_), .Y(_1329_) );
	OAI21X1 OAI21X1_12 ( .A(_1328_), .B(_1140_), .C(_1329_), .Y(_1330_) );
	NOR2X1 NOR2X1_54 ( .A(_1327_), .B(_1330_), .Y(_1331_) );
	NAND3X1 NAND3X1_15 ( .A(_1323_), .B(_1324_), .C(_1331_), .Y(_1332_) );
	INVX1 INVX1_51 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_1333_) );
	NAND2X1 NAND2X1_92 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_1119_), .Y(_1334_) );
	OAI21X1 OAI21X1_13 ( .A(_1333_), .B(_1149_), .C(_1334_), .Y(_1335_) );
	INVX1 INVX1_52 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_1336_) );
	INVX1 INVX1_53 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_1337_) );
	OAI22X1 OAI22X1_10 ( .A(_1336_), .B(_1155_), .C(_1153_), .D(_1337_), .Y(_1338_) );
	NOR2X1 NOR2X1_55 ( .A(_1338_), .B(_1335_), .Y(_1339_) );
	AOI22X1 AOI22X1_46 ( .A(_1239_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_1212_), .Y(_1340_) );
	AND2X2 AND2X2_5 ( .A(_1086_), .B(_1101_), .Y(_1341_) );
	AOI22X1 AOI22X1_47 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_1211_), .C(_1341_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_1342_) );
	NAND3X1 NAND3X1_16 ( .A(_1340_), .B(_1342_), .C(_1339_), .Y(_1343_) );
	NOR3X1 NOR3X1_46 ( .A(_1343_), .B(_1321_), .C(_1332_), .Y(_1344_) );
	INVX1 INVX1_54 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_1345_) );
	NAND2X1 NAND2X1_93 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_1174_), .Y(_1346_) );
	OAI21X1 OAI21X1_14 ( .A(_1176_), .B(_1345_), .C(_1346_), .Y(_1347_) );
	AOI21X1 AOI21X1_8 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_1223_), .C(_1347_), .Y(_1348_) );
	INVX1 INVX1_55 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_1349_) );
	INVX1 INVX1_56 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_1350_) );
	OAI22X1 OAI22X1_11 ( .A(_1350_), .B(_1182_), .C(_1183_), .D(_1349_), .Y(_1351_) );
	INVX1 INVX1_57 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_1352_) );
	NAND2X1 NAND2X1_94 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_1192_), .Y(_1353_) );
	OAI21X1 OAI21X1_15 ( .A(_1093_), .B(_1352_), .C(_1353_), .Y(_1354_) );
	NOR2X1 NOR2X1_56 ( .A(_1354_), .B(_1351_), .Y(_1355_) );
	INVX1 INVX1_58 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_1356_) );
	INVX1 INVX1_59 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_1357_) );
	OAI22X1 OAI22X1_12 ( .A(_1188_), .B(_1357_), .C(_1194_), .D(_1356_), .Y(_1358_) );
	INVX1 INVX1_60 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_1359_) );
	NOR2X1 NOR2X1_57 ( .A(_1359_), .B(_1199_), .Y(_1360_) );
	INVX1 INVX1_61 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_1361_) );
	NOR2X1 NOR2X1_58 ( .A(_1361_), .B(_1200_), .Y(_1362_) );
	NOR3X1 NOR3X1_47 ( .A(_1360_), .B(_1358_), .C(_1362_), .Y(_1363_) );
	NAND3X1 NAND3X1_17 ( .A(_1355_), .B(_1348_), .C(_1363_), .Y(_1364_) );
	AOI22X1 AOI22X1_48 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_1204_), .C(_1205_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_1365_) );
	AOI22X1 AOI22X1_49 ( .A(_1207_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_1208_), .Y(_1366_) );
	NAND2X1 NAND2X1_95 ( .A(_1365_), .B(_1366_), .Y(_1367_) );
	AOI22X1 AOI22X1_50 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_1215_), .C(_1214_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_1368_) );
	AOI22X1 AOI22X1_51 ( .A(_1158_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_1165_), .Y(_1369_) );
	NAND2X1 NAND2X1_96 ( .A(_1368_), .B(_1369_), .Y(_1370_) );
	NOR2X1 NOR2X1_59 ( .A(_1367_), .B(_1370_), .Y(_1371_) );
	AOI22X1 AOI22X1_52 ( .A(_1219_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_1220_), .Y(_1372_) );
	AOI22X1 AOI22X1_53 ( .A(_1121_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_1222_), .Y(_1373_) );
	NAND2X1 NAND2X1_97 ( .A(_1372_), .B(_1373_), .Y(_1374_) );
	AOI22X1 AOI22X1_54 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_1226_), .C(_1227_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_1375_) );
	AOI22X1 AOI22X1_55 ( .A(_1229_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_1230_), .Y(_1376_) );
	NAND2X1 NAND2X1_98 ( .A(_1376_), .B(_1375_), .Y(_1377_) );
	NOR2X1 NOR2X1_60 ( .A(_1374_), .B(_1377_), .Y(_1378_) );
	NAND2X1 NAND2X1_99 ( .A(_1378_), .B(_1371_), .Y(_1379_) );
	AOI22X1 AOI22X1_56 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_1236_), .C(_1137_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_1380_) );
	AOI22X1 AOI22X1_57 ( .A(_1160_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_1238_), .Y(_1381_) );
	NAND2X1 NAND2X1_100 ( .A(_1380_), .B(_1381_), .Y(_1382_) );
	AOI22X1 AOI22X1_58 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_1127_), .C(_1247_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_1383_) );
	NAND2X1 NAND2X1_101 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_1242_), .Y(_1384_) );
	NAND2X1 NAND2X1_102 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_1244_), .Y(_1385_) );
	NAND3X1 NAND3X1_18 ( .A(_1384_), .B(_1385_), .C(_1383_), .Y(_1386_) );
	NOR2X1 NOR2X1_61 ( .A(_1386_), .B(_1382_), .Y(_1387_) );
	AOI22X1 AOI22X1_59 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_1251_), .C(_1252_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_1388_) );
	NAND2X1 NAND2X1_103 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_1254_), .Y(_1389_) );
	NAND2X1 NAND2X1_104 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_1256_), .Y(_1390_) );
	NAND3X1 NAND3X1_19 ( .A(_1389_), .B(_1390_), .C(_1388_), .Y(_1391_) );
	AOI22X1 AOI22X1_60 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_1260_), .C(_1259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_1392_) );
	AOI22X1 AOI22X1_61 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_1263_), .C(_1262_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_1393_) );
	NAND2X1 NAND2X1_105 ( .A(_1392_), .B(_1393_), .Y(_1394_) );
	NOR2X1 NOR2X1_62 ( .A(_1394_), .B(_1391_), .Y(_1395_) );
	NAND2X1 NAND2X1_106 ( .A(_1387_), .B(_1395_), .Y(_1396_) );
	NOR3X1 NOR3X1_48 ( .A(_1379_), .B(_1364_), .C(_1396_), .Y(_1397_) );
	AOI21X1 AOI21X1_9 ( .A(wData[21]), .B(_1273_), .C(_1078_), .Y(_1398_) );
	AOI22X1 AOI22X1_62 ( .A(_1276_), .B(wData[17]), .C(wData[1]), .D(_1304_), .Y(_1399_) );
	AOI22X1 AOI22X1_63 ( .A(_1297_), .B(wData[45]), .C(wData[25]), .D(_1280_), .Y(_1400_) );
	NAND3X1 NAND3X1_20 ( .A(_1398_), .B(_1400_), .C(_1399_), .Y(_1401_) );
	NAND3X1 NAND3X1_21 ( .A(wData[49]), .B(_1274_), .C(_1308_), .Y(_1402_) );
	AOI22X1 AOI22X1_64 ( .A(wData[61]), .B(_1296_), .C(_1284_), .D(wData[5]), .Y(_1403_) );
	AND2X2 AND2X2_6 ( .A(_1403_), .B(_1402_), .Y(_1404_) );
	AOI22X1 AOI22X1_65 ( .A(_1293_), .B(wData[57]), .C(wData[41]), .D(_1300_), .Y(_1405_) );
	AOI22X1 AOI22X1_66 ( .A(wData[53]), .B(_1294_), .C(_1290_), .D(wData[33]), .Y(_1406_) );
	AND2X2 AND2X2_7 ( .A(_1406_), .B(_1405_), .Y(_1407_) );
	AOI22X1 AOI22X1_67 ( .A(_1310_), .B(wData[9]), .C(wData[13]), .D(_1311_), .Y(_1408_) );
	AOI22X1 AOI22X1_68 ( .A(_1286_), .B(wData[29]), .C(wData[37]), .D(_1302_), .Y(_1409_) );
	AND2X2 AND2X2_8 ( .A(_1408_), .B(_1409_), .Y(_1410_) );
	NAND3X1 NAND3X1_22 ( .A(_1404_), .B(_1410_), .C(_1407_), .Y(_1411_) );
	NOR2X1 NOR2X1_63 ( .A(_1401_), .B(_1411_), .Y(_1412_) );
	AOI21X1 AOI21X1_10 ( .A(_1344_), .B(_1397_), .C(_1412_), .Y(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_1_) );
	AOI21X1 AOI21X1_11 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_1317_), .C(_1079_), .Y(_1413_) );
	INVX1 INVX1_62 ( .A(_1176_), .Y(_1414_) );
	AOI22X1 AOI22X1_69 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_1087_), .C(_1414_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_1415_) );
	INVX1 INVX1_63 ( .A(_1188_), .Y(_1416_) );
	AOI22X1 AOI22X1_70 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_1223_), .C(_1416_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_1417_) );
	NAND3X1 NAND3X1_23 ( .A(_1417_), .B(_1413_), .C(_1415_), .Y(_1418_) );
	AOI22X1 AOI22X1_71 ( .A(_1172_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_1322_), .Y(_1419_) );
	AOI22X1 AOI22X1_72 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_1121_), .C(_1094_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_1420_) );
	INVX1 INVX1_64 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_1421_) );
	NAND2X1 NAND2X1_107 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_1211_), .Y(_1422_) );
	OAI21X1 OAI21X1_16 ( .A(_1421_), .B(_1183_), .C(_1422_), .Y(_1423_) );
	INVX1 INVX1_65 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_1424_) );
	NAND2X1 NAND2X1_108 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_1137_), .Y(_1425_) );
	OAI21X1 OAI21X1_17 ( .A(_1424_), .B(_1140_), .C(_1425_), .Y(_1426_) );
	NOR2X1 NOR2X1_64 ( .A(_1423_), .B(_1426_), .Y(_1427_) );
	NAND3X1 NAND3X1_24 ( .A(_1419_), .B(_1420_), .C(_1427_), .Y(_1428_) );
	INVX1 INVX1_66 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_1429_) );
	NAND2X1 NAND2X1_109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_1119_), .Y(_1430_) );
	OAI21X1 OAI21X1_18 ( .A(_1429_), .B(_1149_), .C(_1430_), .Y(_1431_) );
	INVX1 INVX1_67 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_1432_) );
	INVX1 INVX1_68 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_1433_) );
	OAI22X1 OAI22X1_13 ( .A(_1432_), .B(_1155_), .C(_1153_), .D(_1433_), .Y(_1434_) );
	NOR2X1 NOR2X1_65 ( .A(_1434_), .B(_1431_), .Y(_1435_) );
	AOI22X1 AOI22X1_73 ( .A(_1239_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_1212_), .Y(_1436_) );
	AND2X2 AND2X2_9 ( .A(_1111_), .B(_1133_), .Y(_1437_) );
	AOI22X1 AOI22X1_74 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_1437_), .C(_1341_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_1438_) );
	NAND3X1 NAND3X1_25 ( .A(_1436_), .B(_1438_), .C(_1435_), .Y(_1439_) );
	NOR3X1 NOR3X1_49 ( .A(_1439_), .B(_1418_), .C(_1428_), .Y(_1440_) );
	INVX1 INVX1_69 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_1441_) );
	NOR3X1 NOR3X1_50 ( .A(_1441_), .B(_1106_), .C(_1105_), .Y(_1442_) );
	AND2X2 AND2X2_10 ( .A(_1127_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_1443_) );
	AND2X2 AND2X2_11 ( .A(_1247_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_1444_) );
	NOR3X1 NOR3X1_51 ( .A(_1444_), .B(_1443_), .C(_1442_), .Y(_1445_) );
	INVX1 INVX1_70 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_1446_) );
	INVX1 INVX1_71 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_1447_) );
	OAI22X1 OAI22X1_14 ( .A(_1447_), .B(_1182_), .C(_1132_), .D(_1446_), .Y(_1448_) );
	INVX1 INVX1_72 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_1449_) );
	INVX1 INVX1_73 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_1450_) );
	NAND2X1 NAND2X1_110 ( .A(_1123_), .B(_1124_), .Y(_1451_) );
	OAI22X1 OAI22X1_15 ( .A(_1451_), .B(_1450_), .C(_1449_), .D(_1102_), .Y(_1452_) );
	NOR2X1 NOR2X1_66 ( .A(_1448_), .B(_1452_), .Y(_1453_) );
	INVX1 INVX1_74 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_1454_) );
	NOR3X1 NOR3X1_52 ( .A(_1083_), .B(_1100_), .C(_1091_), .Y(_1455_) );
	NAND2X1 NAND2X1_111 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_1455_), .Y(_1456_) );
	OAI21X1 OAI21X1_19 ( .A(_1112_), .B(_1454_), .C(_1456_), .Y(_1457_) );
	INVX1 INVX1_75 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_1458_) );
	INVX1 INVX1_76 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_1459_) );
	OAI22X1 OAI22X1_16 ( .A(_1199_), .B(_1459_), .C(_1458_), .D(_1200_), .Y(_1460_) );
	NOR2X1 NOR2X1_67 ( .A(_1457_), .B(_1460_), .Y(_1461_) );
	NAND3X1 NAND3X1_26 ( .A(_1445_), .B(_1461_), .C(_1453_), .Y(_1462_) );
	AOI22X1 AOI22X1_75 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_1204_), .C(_1205_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_1463_) );
	AOI22X1 AOI22X1_76 ( .A(_1207_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_1208_), .Y(_1464_) );
	NAND2X1 NAND2X1_112 ( .A(_1463_), .B(_1464_), .Y(_1465_) );
	AOI22X1 AOI22X1_77 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_1215_), .C(_1214_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_1466_) );
	AOI22X1 AOI22X1_78 ( .A(_1158_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_1165_), .Y(_1467_) );
	NAND2X1 NAND2X1_113 ( .A(_1466_), .B(_1467_), .Y(_1468_) );
	NOR2X1 NOR2X1_68 ( .A(_1465_), .B(_1468_), .Y(_1469_) );
	AOI22X1 AOI22X1_79 ( .A(_1219_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_1220_), .Y(_1470_) );
	AOI22X1 AOI22X1_80 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_1246_), .C(_1222_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_1471_) );
	NAND2X1 NAND2X1_114 ( .A(_1471_), .B(_1470_), .Y(_1472_) );
	AOI22X1 AOI22X1_81 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_1226_), .C(_1227_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_1473_) );
	AOI22X1 AOI22X1_82 ( .A(_1229_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_1230_), .Y(_1474_) );
	NAND2X1 NAND2X1_115 ( .A(_1474_), .B(_1473_), .Y(_1475_) );
	NOR2X1 NOR2X1_69 ( .A(_1472_), .B(_1475_), .Y(_1476_) );
	NAND2X1 NAND2X1_116 ( .A(_1476_), .B(_1469_), .Y(_1477_) );
	AOI22X1 AOI22X1_83 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_1236_), .C(_1235_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_1478_) );
	AOI22X1 AOI22X1_84 ( .A(_1160_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_1238_), .Y(_1479_) );
	NAND2X1 NAND2X1_117 ( .A(_1478_), .B(_1479_), .Y(_1480_) );
	AOI22X1 AOI22X1_85 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_1244_), .C(_1242_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_1481_) );
	AOI22X1 AOI22X1_86 ( .A(_1174_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_1192_), .Y(_1482_) );
	NAND2X1 NAND2X1_118 ( .A(_1482_), .B(_1481_), .Y(_1483_) );
	NOR2X1 NOR2X1_70 ( .A(_1483_), .B(_1480_), .Y(_1484_) );
	AOI22X1 AOI22X1_87 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_1251_), .C(_1252_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_1485_) );
	NAND2X1 NAND2X1_119 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_1254_), .Y(_1486_) );
	NAND2X1 NAND2X1_120 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_1256_), .Y(_1487_) );
	NAND3X1 NAND3X1_27 ( .A(_1486_), .B(_1487_), .C(_1485_), .Y(_1488_) );
	AOI22X1 AOI22X1_88 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_1260_), .C(_1259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_1489_) );
	AOI22X1 AOI22X1_89 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_1263_), .C(_1262_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_1490_) );
	NAND2X1 NAND2X1_121 ( .A(_1489_), .B(_1490_), .Y(_1491_) );
	NOR2X1 NOR2X1_71 ( .A(_1491_), .B(_1488_), .Y(_1492_) );
	NAND2X1 NAND2X1_122 ( .A(_1484_), .B(_1492_), .Y(_1493_) );
	NOR3X1 NOR3X1_53 ( .A(_1477_), .B(_1462_), .C(_1493_), .Y(_1494_) );
	AOI22X1 AOI22X1_90 ( .A(_1300_), .B(wData[42]), .C(wData[38]), .D(_1302_), .Y(_1495_) );
	AOI22X1 AOI22X1_91 ( .A(_1297_), .B(wData[46]), .C(_1304_), .D(wData[2]), .Y(_1496_) );
	NAND2X1 NAND2X1_123 ( .A(_1495_), .B(_1496_), .Y(_1497_) );
	AOI21X1 AOI21X1_12 ( .A(wData[34]), .B(_1290_), .C(_1497_), .Y(_1498_) );
	INVX1 INVX1_77 ( .A(wData[50]), .Y(_1499_) );
	AOI22X1 AOI22X1_92 ( .A(_1310_), .B(wData[10]), .C(wData[14]), .D(_1311_), .Y(_1500_) );
	OAI21X1 OAI21X1_20 ( .A(_1499_), .B(_1309_), .C(_1500_), .Y(_1501_) );
	AOI22X1 AOI22X1_93 ( .A(_1273_), .B(wData[22]), .C(wData[18]), .D(_1276_), .Y(_1502_) );
	NAND2X1 NAND2X1_124 ( .A(wData[26]), .B(_1280_), .Y(_1503_) );
	AOI22X1 AOI22X1_94 ( .A(_1286_), .B(wData[30]), .C(wData[6]), .D(_1284_), .Y(_1504_) );
	NAND3X1 NAND3X1_28 ( .A(_1503_), .B(_1504_), .C(_1502_), .Y(_1505_) );
	NOR2X1 NOR2X1_72 ( .A(_1501_), .B(_1505_), .Y(_1506_) );
	NAND2X1 NAND2X1_125 ( .A(wData[58]), .B(_1293_), .Y(_1507_) );
	NAND2X1 NAND2X1_126 ( .A(wData[54]), .B(_1294_), .Y(_1508_) );
	NAND2X1 NAND2X1_127 ( .A(_1507_), .B(_1508_), .Y(_1509_) );
	AOI21X1 AOI21X1_13 ( .A(wData[62]), .B(_1296_), .C(_1509_), .Y(_1510_) );
	NAND3X1 NAND3X1_29 ( .A(_1498_), .B(_1510_), .C(_1506_), .Y(_1511_) );
	NOR2X1 NOR2X1_73 ( .A(_1078_), .B(_1511_), .Y(_1512_) );
	AOI21X1 AOI21X1_14 ( .A(_1440_), .B(_1494_), .C(_1512_), .Y(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_2_) );
	AOI21X1 AOI21X1_15 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_1322_), .C(_1079_), .Y(_1513_) );
	AOI22X1 AOI22X1_95 ( .A(_1094_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_1414_), .Y(_1514_) );
	AOI22X1 AOI22X1_96 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_1416_), .C(_1172_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_1515_) );
	NAND3X1 NAND3X1_30 ( .A(_1515_), .B(_1513_), .C(_1514_), .Y(_1516_) );
	AOI22X1 AOI22X1_97 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_1121_), .C(_1119_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_1517_) );
	AOI22X1 AOI22X1_98 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_1192_), .C(_1317_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_1518_) );
	INVX1 INVX1_78 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_1519_) );
	INVX1 INVX1_79 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_1520_) );
	OAI22X1 OAI22X1_17 ( .A(_1519_), .B(_1134_), .C(_1183_), .D(_1520_), .Y(_1521_) );
	INVX1 INVX1_80 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_1522_) );
	NAND2X1 NAND2X1_128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_1235_), .Y(_1523_) );
	OAI21X1 OAI21X1_21 ( .A(_1522_), .B(_1140_), .C(_1523_), .Y(_1524_) );
	NOR2X1 NOR2X1_74 ( .A(_1521_), .B(_1524_), .Y(_1525_) );
	NAND3X1 NAND3X1_31 ( .A(_1517_), .B(_1518_), .C(_1525_), .Y(_1526_) );
	AND2X2 AND2X2_12 ( .A(_1148_), .B(_1082_), .Y(_1527_) );
	AOI22X1 AOI22X1_99 ( .A(_1087_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_1527_), .Y(_1528_) );
	AND2X2 AND2X2_13 ( .A(_1146_), .B(_1111_), .Y(_1529_) );
	AND2X2 AND2X2_14 ( .A(_1154_), .B(_1111_), .Y(_1530_) );
	AOI22X1 AOI22X1_100 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_1530_), .C(_1529_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_1531_) );
	NAND2X1 NAND2X1_129 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_1239_), .Y(_1532_) );
	NAND2X1 NAND2X1_130 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_1212_), .Y(_1533_) );
	NAND2X1 NAND2X1_131 ( .A(_1532_), .B(_1533_), .Y(_1534_) );
	INVX1 INVX1_81 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_1535_) );
	NAND2X1 NAND2X1_132 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_1211_), .Y(_1536_) );
	OAI21X1 OAI21X1_22 ( .A(_1535_), .B(_1164_), .C(_1536_), .Y(_1537_) );
	NOR2X1 NOR2X1_75 ( .A(_1534_), .B(_1537_), .Y(_1538_) );
	NAND3X1 NAND3X1_32 ( .A(_1528_), .B(_1531_), .C(_1538_), .Y(_1539_) );
	NOR3X1 NOR3X1_54 ( .A(_1526_), .B(_1516_), .C(_1539_), .Y(_1540_) );
	INVX1 INVX1_82 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_1541_) );
	NAND2X1 NAND2X1_133 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_1127_), .Y(_1542_) );
	OAI21X1 OAI21X1_23 ( .A(_1132_), .B(_1541_), .C(_1542_), .Y(_1543_) );
	AOI21X1 AOI21X1_16 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_1107_), .C(_1543_), .Y(_1544_) );
	INVX1 INVX1_83 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_1545_) );
	INVX1 INVX1_84 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_1546_) );
	OAI22X1 OAI22X1_18 ( .A(_1451_), .B(_1546_), .C(_1545_), .D(_1102_), .Y(_1547_) );
	INVX1 INVX1_85 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_1548_) );
	NAND2X1 NAND2X1_134 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_1247_), .Y(_1549_) );
	OAI21X1 OAI21X1_24 ( .A(_1112_), .B(_1548_), .C(_1549_), .Y(_1550_) );
	NOR2X1 NOR2X1_76 ( .A(_1550_), .B(_1547_), .Y(_1551_) );
	INVX1 INVX1_86 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_1552_) );
	INVX1 INVX1_87 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_1553_) );
	OAI22X1 OAI22X1_19 ( .A(_1199_), .B(_1553_), .C(_1552_), .D(_1200_), .Y(_1554_) );
	INVX1 INVX1_88 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_1555_) );
	NAND2X1 NAND2X1_135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_1246_), .Y(_1556_) );
	OAI21X1 OAI21X1_25 ( .A(_1555_), .B(_1182_), .C(_1556_), .Y(_1557_) );
	NOR2X1 NOR2X1_77 ( .A(_1557_), .B(_1554_), .Y(_1558_) );
	NAND3X1 NAND3X1_33 ( .A(_1544_), .B(_1558_), .C(_1551_), .Y(_1559_) );
	AOI22X1 AOI22X1_101 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_1204_), .C(_1205_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_1560_) );
	AOI22X1 AOI22X1_102 ( .A(_1207_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_1208_), .Y(_1561_) );
	NAND2X1 NAND2X1_136 ( .A(_1560_), .B(_1561_), .Y(_1562_) );
	AOI22X1 AOI22X1_103 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_1215_), .C(_1214_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_1563_) );
	AOI22X1 AOI22X1_104 ( .A(_1158_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_1165_), .Y(_1564_) );
	NAND2X1 NAND2X1_137 ( .A(_1563_), .B(_1564_), .Y(_1565_) );
	NOR2X1 NOR2X1_78 ( .A(_1562_), .B(_1565_), .Y(_1566_) );
	AOI22X1 AOI22X1_105 ( .A(_1219_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_1220_), .Y(_1567_) );
	AOI22X1 AOI22X1_106 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_1455_), .C(_1222_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_1568_) );
	NAND2X1 NAND2X1_138 ( .A(_1568_), .B(_1567_), .Y(_1569_) );
	AOI22X1 AOI22X1_107 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_1226_), .C(_1227_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_1570_) );
	AOI22X1 AOI22X1_108 ( .A(_1229_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_1230_), .Y(_1571_) );
	NAND2X1 NAND2X1_139 ( .A(_1571_), .B(_1570_), .Y(_1572_) );
	NOR2X1 NOR2X1_79 ( .A(_1569_), .B(_1572_), .Y(_1573_) );
	NAND2X1 NAND2X1_140 ( .A(_1573_), .B(_1566_), .Y(_1574_) );
	AOI22X1 AOI22X1_109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_1236_), .C(_1137_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_1575_) );
	AOI22X1 AOI22X1_110 ( .A(_1160_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_1238_), .Y(_1576_) );
	NAND2X1 NAND2X1_141 ( .A(_1575_), .B(_1576_), .Y(_1577_) );
	AOI22X1 AOI22X1_111 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_1244_), .C(_1242_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_1578_) );
	AOI22X1 AOI22X1_112 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_1174_), .C(_1223_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_1579_) );
	NAND2X1 NAND2X1_142 ( .A(_1579_), .B(_1578_), .Y(_1580_) );
	NOR2X1 NOR2X1_80 ( .A(_1580_), .B(_1577_), .Y(_1581_) );
	AOI22X1 AOI22X1_113 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_1251_), .C(_1252_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_1582_) );
	NAND2X1 NAND2X1_143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_1254_), .Y(_1583_) );
	NAND2X1 NAND2X1_144 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_1256_), .Y(_1584_) );
	NAND3X1 NAND3X1_34 ( .A(_1583_), .B(_1584_), .C(_1582_), .Y(_1585_) );
	AOI22X1 AOI22X1_114 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_1260_), .C(_1259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_1586_) );
	AOI22X1 AOI22X1_115 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_1263_), .C(_1262_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_1587_) );
	NAND2X1 NAND2X1_145 ( .A(_1586_), .B(_1587_), .Y(_1588_) );
	NOR2X1 NOR2X1_81 ( .A(_1588_), .B(_1585_), .Y(_1589_) );
	NAND2X1 NAND2X1_146 ( .A(_1581_), .B(_1589_), .Y(_1590_) );
	NOR3X1 NOR3X1_55 ( .A(_1574_), .B(_1559_), .C(_1590_), .Y(_1591_) );
	NAND2X1 NAND2X1_147 ( .A(wData[59]), .B(_1293_), .Y(_1592_) );
	OAI21X1 OAI21X1_26 ( .A(_1077_), .B(wBusy_bF_buf2), .C(_1592_), .Y(_1593_) );
	NAND2X1 NAND2X1_148 ( .A(wData[7]), .B(_1284_), .Y(_1594_) );
	NAND2X1 NAND2X1_149 ( .A(wData[55]), .B(_1294_), .Y(_1595_) );
	AOI22X1 AOI22X1_116 ( .A(wData[63]), .B(_1296_), .C(_1286_), .D(wData[31]), .Y(_1596_) );
	NAND3X1 NAND3X1_35 ( .A(_1594_), .B(_1595_), .C(_1596_), .Y(_1597_) );
	OR2X2 OR2X2_8 ( .A(_1597_), .B(_1593_), .Y(_1598_) );
	INVX1 INVX1_89 ( .A(wData[51]), .Y(_1599_) );
	NAND2X1 NAND2X1_150 ( .A(wData[47]), .B(_1297_), .Y(_1600_) );
	OAI21X1 OAI21X1_27 ( .A(_1599_), .B(_1309_), .C(_1600_), .Y(_1601_) );
	AOI21X1 AOI21X1_17 ( .A(wData[3]), .B(_1304_), .C(_1601_), .Y(_1602_) );
	AOI22X1 AOI22X1_117 ( .A(_1310_), .B(wData[11]), .C(wData[15]), .D(_1311_), .Y(_1603_) );
	AOI22X1 AOI22X1_118 ( .A(_1273_), .B(wData[23]), .C(wData[27]), .D(_1280_), .Y(_1604_) );
	AND2X2 AND2X2_15 ( .A(_1603_), .B(_1604_), .Y(_1605_) );
	NAND2X1 NAND2X1_151 ( .A(wData[39]), .B(_1302_), .Y(_1606_) );
	NAND2X1 NAND2X1_152 ( .A(wData[43]), .B(_1300_), .Y(_1607_) );
	NAND2X1 NAND2X1_153 ( .A(_1606_), .B(_1607_), .Y(_1608_) );
	NAND2X1 NAND2X1_154 ( .A(wData[19]), .B(_1276_), .Y(_1609_) );
	NAND2X1 NAND2X1_155 ( .A(wData[35]), .B(_1290_), .Y(_1610_) );
	NAND2X1 NAND2X1_156 ( .A(_1609_), .B(_1610_), .Y(_1611_) );
	NOR2X1 NOR2X1_82 ( .A(_1608_), .B(_1611_), .Y(_1612_) );
	NAND3X1 NAND3X1_36 ( .A(_1605_), .B(_1602_), .C(_1612_), .Y(_1613_) );
	NOR2X1 NOR2X1_83 ( .A(_1598_), .B(_1613_), .Y(_1614_) );
	AOI21X1 AOI21X1_18 ( .A(_1540_), .B(_1591_), .C(_1614_), .Y(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_3_) );
	INVX1 INVX1_90 ( .A(wSelec[33]), .Y(_1615_) );
	NOR2X1 NOR2X1_84 ( .A(wBusy_bF_buf1), .B(_1615_), .Y(_1616_) );
	INVX1 INVX1_91 ( .A(_1616_), .Y(_1617_) );
	INVX1 INVX1_92 ( .A(wSelec[43]), .Y(_1618_) );
	NAND2X1 NAND2X1_157 ( .A(wSelec[42]), .B(_1618_), .Y(_1619_) );
	INVX2 INVX2_3 ( .A(_1619_), .Y(_1620_) );
	OR2X2 OR2X2_9 ( .A(wSelec[39]), .B(wSelec[38]), .Y(_1621_) );
	INVX1 INVX1_93 ( .A(wSelec[41]), .Y(_1622_) );
	NAND2X1 NAND2X1_158 ( .A(wSelec[40]), .B(_1622_), .Y(_1623_) );
	NOR2X1 NOR2X1_85 ( .A(_1621_), .B(_1623_), .Y(_1624_) );
	AND2X2 AND2X2_16 ( .A(_1624_), .B(_1620_), .Y(_1625_) );
	AOI21X1 AOI21X1_19 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_1625_), .C(_1617_), .Y(_1626_) );
	INVX1 INVX1_94 ( .A(wSelec[39]), .Y(_1627_) );
	NAND2X1 NAND2X1_159 ( .A(wSelec[38]), .B(_1627_), .Y(_1628_) );
	OR2X2 OR2X2_10 ( .A(wSelec[40]), .B(wSelec[41]), .Y(_1629_) );
	NOR2X1 NOR2X1_86 ( .A(_1629_), .B(_1628_), .Y(_1630_) );
	NAND2X1 NAND2X1_160 ( .A(_1620_), .B(_1630_), .Y(_1631_) );
	INVX1 INVX1_95 ( .A(_1631_), .Y(_1632_) );
	INVX1 INVX1_96 ( .A(wSelec[38]), .Y(_1633_) );
	NAND2X1 NAND2X1_161 ( .A(wSelec[39]), .B(_1633_), .Y(_1634_) );
	INVX1 INVX1_97 ( .A(wSelec[40]), .Y(_1635_) );
	NAND2X1 NAND2X1_162 ( .A(wSelec[41]), .B(_1635_), .Y(_1636_) );
	NOR2X1 NOR2X1_87 ( .A(_1634_), .B(_1636_), .Y(_1637_) );
	NAND2X1 NAND2X1_163 ( .A(wSelec[42]), .B(wSelec[43]), .Y(_1638_) );
	INVX1 INVX1_98 ( .A(_1638_), .Y(_1639_) );
	NAND2X1 NAND2X1_164 ( .A(_1639_), .B(_1637_), .Y(_1640_) );
	INVX1 INVX1_99 ( .A(_1640_), .Y(_1641_) );
	AOI22X1 AOI22X1_119 ( .A(_1632_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_1641_), .Y(_1642_) );
	OR2X2 OR2X2_11 ( .A(_1628_), .B(_1629_), .Y(_1643_) );
	OR2X2 OR2X2_12 ( .A(wSelec[42]), .B(wSelec[43]), .Y(_1644_) );
	NOR2X1 NOR2X1_88 ( .A(_1644_), .B(_1643_), .Y(_1645_) );
	NOR2X1 NOR2X1_89 ( .A(_1623_), .B(_1628_), .Y(_1646_) );
	INVX1 INVX1_100 ( .A(wSelec[42]), .Y(_1647_) );
	NAND2X1 NAND2X1_165 ( .A(wSelec[43]), .B(_1647_), .Y(_1648_) );
	INVX2 INVX2_4 ( .A(_1648_), .Y(_1649_) );
	NAND2X1 NAND2X1_166 ( .A(_1649_), .B(_1646_), .Y(_1650_) );
	INVX1 INVX1_101 ( .A(_1650_), .Y(_1651_) );
	AOI22X1 AOI22X1_120 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_1645_), .C(_1651_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_1652_) );
	NAND3X1 NAND3X1_37 ( .A(_1626_), .B(_1652_), .C(_1642_), .Y(_1653_) );
	NOR2X1 NOR2X1_90 ( .A(wSelec[39]), .B(wSelec[38]), .Y(_1654_) );
	NOR2X1 NOR2X1_91 ( .A(wSelec[40]), .B(wSelec[41]), .Y(_1655_) );
	NAND2X1 NAND2X1_167 ( .A(_1654_), .B(_1655_), .Y(_1656_) );
	NOR2X1 NOR2X1_92 ( .A(_1619_), .B(_1656_), .Y(_1657_) );
	NAND2X1 NAND2X1_168 ( .A(wSelec[39]), .B(wSelec[38]), .Y(_1658_) );
	NOR3X1 NOR3X1_56 ( .A(_1629_), .B(_1658_), .C(_1619_), .Y(_1659_) );
	AOI22X1 AOI22X1_121 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_1659_), .C(_1657_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_1660_) );
	INVX1 INVX1_102 ( .A(_1644_), .Y(_1661_) );
	NOR2X1 NOR2X1_93 ( .A(_1629_), .B(_1634_), .Y(_1662_) );
	AND2X2 AND2X2_17 ( .A(_1662_), .B(_1661_), .Y(_1663_) );
	NAND2X1 NAND2X1_169 ( .A(wSelec[40]), .B(wSelec[41]), .Y(_1664_) );
	NOR3X1 NOR3X1_57 ( .A(_1638_), .B(_1658_), .C(_1664_), .Y(_1665_) );
	AOI22X1 AOI22X1_122 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_1665_), .C(_1663_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_1666_) );
	INVX1 INVX1_103 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_1667_) );
	INVX1 INVX1_104 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_1668_) );
	NOR2X1 NOR2X1_94 ( .A(_1628_), .B(_1636_), .Y(_1669_) );
	NAND2X1 NAND2X1_170 ( .A(_1639_), .B(_1669_), .Y(_1670_) );
	NOR2X1 NOR2X1_95 ( .A(_1658_), .B(_1664_), .Y(_1671_) );
	NAND2X1 NAND2X1_171 ( .A(_1671_), .B(_1649_), .Y(_1672_) );
	OAI22X1 OAI22X1_20 ( .A(_1667_), .B(_1672_), .C(_1670_), .D(_1668_), .Y(_1673_) );
	INVX1 INVX1_105 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_1674_) );
	NOR3X1 NOR3X1_58 ( .A(_1619_), .B(_1634_), .C(_1636_), .Y(_1675_) );
	NAND2X1 NAND2X1_172 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_1675_), .Y(_1676_) );
	NOR2X1 NOR2X1_96 ( .A(_1658_), .B(_1623_), .Y(_1677_) );
	NAND2X1 NAND2X1_173 ( .A(_1649_), .B(_1677_), .Y(_1678_) );
	OAI21X1 OAI21X1_28 ( .A(_1674_), .B(_1678_), .C(_1676_), .Y(_1679_) );
	NOR2X1 NOR2X1_97 ( .A(_1673_), .B(_1679_), .Y(_1680_) );
	NAND3X1 NAND3X1_38 ( .A(_1660_), .B(_1666_), .C(_1680_), .Y(_1681_) );
	INVX1 INVX1_106 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_1682_) );
	INVX1 INVX1_107 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_1683_) );
	NOR2X1 NOR2X1_98 ( .A(_1623_), .B(_1634_), .Y(_1684_) );
	NAND2X1 NAND2X1_174 ( .A(_1620_), .B(_1684_), .Y(_1685_) );
	NOR2X1 NOR2X1_99 ( .A(_1621_), .B(_1636_), .Y(_1686_) );
	NAND2X1 NAND2X1_175 ( .A(_1620_), .B(_1686_), .Y(_1687_) );
	OAI22X1 OAI22X1_21 ( .A(_1687_), .B(_1682_), .C(_1683_), .D(_1685_), .Y(_1688_) );
	INVX1 INVX1_108 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_1689_) );
	INVX1 INVX1_109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_1690_) );
	NAND2X1 NAND2X1_176 ( .A(_1649_), .B(_1684_), .Y(_1691_) );
	NOR2X1 NOR2X1_100 ( .A(_1658_), .B(_1629_), .Y(_1692_) );
	NAND2X1 NAND2X1_177 ( .A(_1649_), .B(_1692_), .Y(_1693_) );
	OAI22X1 OAI22X1_22 ( .A(_1689_), .B(_1693_), .C(_1691_), .D(_1690_), .Y(_1694_) );
	NOR2X1 NOR2X1_101 ( .A(_1694_), .B(_1688_), .Y(_1695_) );
	NOR3X1 NOR3X1_59 ( .A(_1628_), .B(_1664_), .C(_1648_), .Y(_1696_) );
	NAND2X1 NAND2X1_178 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_1696_), .Y(_1697_) );
	NOR3X1 NOR3X1_60 ( .A(_1636_), .B(_1658_), .C(_1648_), .Y(_1698_) );
	NAND2X1 NAND2X1_179 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_1698_), .Y(_1699_) );
	NAND2X1 NAND2X1_180 ( .A(_1697_), .B(_1699_), .Y(_1700_) );
	INVX1 INVX1_110 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_1701_) );
	NAND2X1 NAND2X1_181 ( .A(_1639_), .B(_1624_), .Y(_1702_) );
	NOR3X1 NOR3X1_61 ( .A(_1634_), .B(_1636_), .C(_1648_), .Y(_1703_) );
	NAND2X1 NAND2X1_182 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_1703_), .Y(_1704_) );
	OAI21X1 OAI21X1_29 ( .A(_1701_), .B(_1702_), .C(_1704_), .Y(_1705_) );
	NOR2X1 NOR2X1_102 ( .A(_1700_), .B(_1705_), .Y(_1706_) );
	NAND2X1 NAND2X1_183 ( .A(_1695_), .B(_1706_), .Y(_1707_) );
	NOR3X1 NOR3X1_62 ( .A(_1653_), .B(_1707_), .C(_1681_), .Y(_1708_) );
	NAND2X1 NAND2X1_184 ( .A(_1620_), .B(_1677_), .Y(_1709_) );
	INVX1 INVX1_111 ( .A(_1709_), .Y(_1710_) );
	INVX1 INVX1_112 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_1711_) );
	NOR3X1 NOR3X1_63 ( .A(_1621_), .B(_1644_), .C(_1623_), .Y(_1712_) );
	NAND2X1 NAND2X1_185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_1712_), .Y(_1713_) );
	NAND2X1 NAND2X1_186 ( .A(_1661_), .B(_1684_), .Y(_1714_) );
	OAI21X1 OAI21X1_30 ( .A(_1714_), .B(_1711_), .C(_1713_), .Y(_1715_) );
	AOI21X1 AOI21X1_20 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_1710_), .C(_1715_), .Y(_1716_) );
	INVX1 INVX1_113 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_1717_) );
	INVX1 INVX1_114 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_1718_) );
	NOR2X1 NOR2X1_103 ( .A(_1664_), .B(_1621_), .Y(_1719_) );
	NAND2X1 NAND2X1_187 ( .A(_1620_), .B(_1719_), .Y(_1720_) );
	NAND2X1 NAND2X1_188 ( .A(_1661_), .B(_1646_), .Y(_1721_) );
	OAI22X1 OAI22X1_23 ( .A(_1718_), .B(_1720_), .C(_1721_), .D(_1717_), .Y(_1722_) );
	INVX1 INVX1_115 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_1723_) );
	INVX1 INVX1_116 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_1724_) );
	NAND2X1 NAND2X1_189 ( .A(_1620_), .B(_1646_), .Y(_1725_) );
	NAND2X1 NAND2X1_190 ( .A(_1661_), .B(_1692_), .Y(_1726_) );
	OAI22X1 OAI22X1_24 ( .A(_1723_), .B(_1726_), .C(_1725_), .D(_1724_), .Y(_1727_) );
	NOR2X1 NOR2X1_104 ( .A(_1722_), .B(_1727_), .Y(_1728_) );
	INVX1 INVX1_117 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_1729_) );
	NOR3X1 NOR3X1_64 ( .A(_1644_), .B(_1658_), .C(_1623_), .Y(_1730_) );
	NAND2X1 NAND2X1_191 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_1730_), .Y(_1731_) );
	OR2X2 OR2X2_13 ( .A(_1656_), .B(_1638_), .Y(_1732_) );
	OAI21X1 OAI21X1_31 ( .A(_1729_), .B(_1732_), .C(_1731_), .Y(_1733_) );
	INVX1 INVX1_118 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_1734_) );
	INVX1 INVX1_119 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_1735_) );
	NOR2X1 NOR2X1_105 ( .A(_1664_), .B(_1634_), .Y(_1736_) );
	NAND2X1 NAND2X1_192 ( .A(_1620_), .B(_1736_), .Y(_1737_) );
	NAND2X1 NAND2X1_193 ( .A(_1639_), .B(_1630_), .Y(_1738_) );
	OAI22X1 OAI22X1_25 ( .A(_1737_), .B(_1735_), .C(_1734_), .D(_1738_), .Y(_1739_) );
	NOR2X1 NOR2X1_106 ( .A(_1733_), .B(_1739_), .Y(_1740_) );
	NAND3X1 NAND3X1_39 ( .A(_1716_), .B(_1740_), .C(_1728_), .Y(_1741_) );
	NOR3X1 NOR3X1_65 ( .A(_1621_), .B(_1629_), .C(_1644_), .Y(_1742_) );
	NOR3X1 NOR3X1_66 ( .A(_1638_), .B(_1664_), .C(_1628_), .Y(_1743_) );
	AOI22X1 AOI22X1_123 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_1742_), .C(_1743_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_1744_) );
	NOR3X1 NOR3X1_67 ( .A(_1638_), .B(_1664_), .C(_1634_), .Y(_1745_) );
	NOR3X1 NOR3X1_68 ( .A(_1638_), .B(_1658_), .C(_1636_), .Y(_1746_) );
	AOI22X1 AOI22X1_124 ( .A(_1745_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_1746_), .Y(_1747_) );
	NAND2X1 NAND2X1_194 ( .A(_1744_), .B(_1747_), .Y(_1748_) );
	NOR3X1 NOR3X1_69 ( .A(_1636_), .B(_1621_), .C(_1648_), .Y(_1749_) );
	NOR3X1 NOR3X1_70 ( .A(_1628_), .B(_1636_), .C(_1648_), .Y(_1750_) );
	AOI22X1 AOI22X1_125 ( .A(_1749_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_1750_), .Y(_1751_) );
	NOR3X1 NOR3X1_71 ( .A(_1619_), .B(_1664_), .C(_1628_), .Y(_1752_) );
	NOR3X1 NOR3X1_72 ( .A(_1658_), .B(_1664_), .C(_1619_), .Y(_1753_) );
	AOI22X1 AOI22X1_126 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_1753_), .C(_1752_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_1754_) );
	NAND2X1 NAND2X1_195 ( .A(_1754_), .B(_1751_), .Y(_1755_) );
	NOR2X1 NOR2X1_107 ( .A(_1748_), .B(_1755_), .Y(_1756_) );
	NOR3X1 NOR3X1_73 ( .A(_1644_), .B(_1664_), .C(_1628_), .Y(_1757_) );
	NOR3X1 NOR3X1_74 ( .A(_1644_), .B(_1664_), .C(_1634_), .Y(_1758_) );
	AOI22X1 AOI22X1_127 ( .A(_1757_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_1758_), .Y(_1759_) );
	NOR3X1 NOR3X1_75 ( .A(_1644_), .B(_1658_), .C(_1636_), .Y(_1760_) );
	NOR3X1 NOR3X1_76 ( .A(_1619_), .B(_1629_), .C(_1634_), .Y(_1761_) );
	AOI22X1 AOI22X1_128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_1760_), .C(_1761_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_1762_) );
	NAND2X1 NAND2X1_196 ( .A(_1759_), .B(_1762_), .Y(_1763_) );
	NOR3X1 NOR3X1_77 ( .A(_1658_), .B(_1664_), .C(_1644_), .Y(_1764_) );
	NOR3X1 NOR3X1_78 ( .A(_1634_), .B(_1629_), .C(_1648_), .Y(_1765_) );
	AOI22X1 AOI22X1_129 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_1764_), .C(_1765_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_1766_) );
	NOR3X1 NOR3X1_79 ( .A(_1621_), .B(_1629_), .C(_1648_), .Y(_1767_) );
	NOR3X1 NOR3X1_80 ( .A(_1621_), .B(_1664_), .C(_1648_), .Y(_1768_) );
	AOI22X1 AOI22X1_130 ( .A(_1767_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_1768_), .Y(_1769_) );
	NAND2X1 NAND2X1_197 ( .A(_1769_), .B(_1766_), .Y(_1770_) );
	NOR2X1 NOR2X1_108 ( .A(_1763_), .B(_1770_), .Y(_1771_) );
	NAND2X1 NAND2X1_198 ( .A(_1771_), .B(_1756_), .Y(_1772_) );
	NOR3X1 NOR3X1_81 ( .A(_1619_), .B(_1658_), .C(_1636_), .Y(_1773_) );
	NOR3X1 NOR3X1_82 ( .A(_1629_), .B(_1638_), .C(_1634_), .Y(_1774_) );
	AOI22X1 AOI22X1_131 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_1774_), .C(_1773_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_1775_) );
	NOR3X1 NOR3X1_83 ( .A(_1623_), .B(_1621_), .C(_1648_), .Y(_1776_) );
	NOR3X1 NOR3X1_84 ( .A(_1634_), .B(_1664_), .C(_1648_), .Y(_1777_) );
	AOI22X1 AOI22X1_132 ( .A(_1776_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_1777_), .Y(_1778_) );
	NAND2X1 NAND2X1_199 ( .A(_1775_), .B(_1778_), .Y(_1779_) );
	NOR3X1 NOR3X1_85 ( .A(_1619_), .B(_1628_), .C(_1636_), .Y(_1780_) );
	NAND2X1 NAND2X1_200 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_1780_), .Y(_1781_) );
	NOR3X1 NOR3X1_86 ( .A(_1638_), .B(_1658_), .C(_1623_), .Y(_1782_) );
	NAND2X1 NAND2X1_201 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_1782_), .Y(_1783_) );
	NOR3X1 NOR3X1_87 ( .A(_1621_), .B(_1664_), .C(_1644_), .Y(_1784_) );
	NOR3X1 NOR3X1_88 ( .A(_1621_), .B(_1638_), .C(_1636_), .Y(_1785_) );
	AOI22X1 AOI22X1_133 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_1784_), .C(_1785_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_1786_) );
	NAND3X1 NAND3X1_40 ( .A(_1781_), .B(_1783_), .C(_1786_), .Y(_1787_) );
	NOR2X1 NOR2X1_109 ( .A(_1787_), .B(_1779_), .Y(_1788_) );
	NOR3X1 NOR3X1_89 ( .A(_1621_), .B(_1644_), .C(_1636_), .Y(_1789_) );
	NOR3X1 NOR3X1_90 ( .A(_1623_), .B(_1638_), .C(_1628_), .Y(_1790_) );
	AOI22X1 AOI22X1_134 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_1789_), .C(_1790_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_1791_) );
	NOR3X1 NOR3X1_91 ( .A(_1623_), .B(_1638_), .C(_1634_), .Y(_1792_) );
	NAND2X1 NAND2X1_202 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_1792_), .Y(_1793_) );
	NOR3X1 NOR3X1_92 ( .A(_1628_), .B(_1629_), .C(_1648_), .Y(_1794_) );
	NAND2X1 NAND2X1_203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_1794_), .Y(_1795_) );
	NAND3X1 NAND3X1_41 ( .A(_1793_), .B(_1795_), .C(_1791_), .Y(_1796_) );
	NOR3X1 NOR3X1_93 ( .A(_1628_), .B(_1644_), .C(_1636_), .Y(_1797_) );
	NOR3X1 NOR3X1_94 ( .A(_1638_), .B(_1664_), .C(_1621_), .Y(_1798_) );
	AOI22X1 AOI22X1_135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_1798_), .C(_1797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_1799_) );
	NOR3X1 NOR3X1_95 ( .A(_1634_), .B(_1644_), .C(_1636_), .Y(_1800_) );
	NOR3X1 NOR3X1_96 ( .A(_1638_), .B(_1658_), .C(_1629_), .Y(_1801_) );
	AOI22X1 AOI22X1_136 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_1801_), .C(_1800_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_1802_) );
	NAND2X1 NAND2X1_204 ( .A(_1799_), .B(_1802_), .Y(_1803_) );
	NOR2X1 NOR2X1_110 ( .A(_1803_), .B(_1796_), .Y(_1804_) );
	NAND2X1 NAND2X1_205 ( .A(_1788_), .B(_1804_), .Y(_1805_) );
	NOR3X1 NOR3X1_97 ( .A(_1772_), .B(_1741_), .C(_1805_), .Y(_1806_) );
	INVX1 INVX1_120 ( .A(wSelec[35]), .Y(_1807_) );
	NAND2X1 NAND2X1_206 ( .A(wSelec[34]), .B(_1807_), .Y(_1808_) );
	INVX1 INVX1_121 ( .A(wSelec[37]), .Y(_1809_) );
	NAND2X1 NAND2X1_207 ( .A(wSelec[36]), .B(_1809_), .Y(_1810_) );
	NOR2X1 NOR2X1_111 ( .A(_1808_), .B(_1810_), .Y(_1811_) );
	NOR2X1 NOR2X1_112 ( .A(wSelec[35]), .B(wSelec[34]), .Y(_1812_) );
	INVX1 INVX1_122 ( .A(_1812_), .Y(_1813_) );
	NOR2X1 NOR2X1_113 ( .A(_1810_), .B(_1813_), .Y(_1814_) );
	AOI22X1 AOI22X1_137 ( .A(wData[20]), .B(_1811_), .C(_1814_), .D(wData[16]), .Y(_1815_) );
	INVX1 INVX1_123 ( .A(wSelec[34]), .Y(_1816_) );
	NAND2X1 NAND2X1_208 ( .A(wSelec[35]), .B(_1816_), .Y(_1817_) );
	NOR2X1 NOR2X1_114 ( .A(_1817_), .B(_1810_), .Y(_1818_) );
	NAND2X1 NAND2X1_209 ( .A(wData[24]), .B(_1818_), .Y(_1819_) );
	INVX1 INVX1_124 ( .A(wSelec[36]), .Y(_1820_) );
	NAND2X1 NAND2X1_210 ( .A(_1820_), .B(_1809_), .Y(_1821_) );
	NOR2X1 NOR2X1_115 ( .A(_1808_), .B(_1821_), .Y(_1822_) );
	NAND2X1 NAND2X1_211 ( .A(wSelec[35]), .B(wSelec[34]), .Y(_1823_) );
	NOR2X1 NOR2X1_116 ( .A(_1823_), .B(_1810_), .Y(_1824_) );
	AOI22X1 AOI22X1_138 ( .A(_1824_), .B(wData[28]), .C(wData[4]), .D(_1822_), .Y(_1825_) );
	NAND3X1 NAND3X1_42 ( .A(_1819_), .B(_1825_), .C(_1815_), .Y(_1826_) );
	NAND2X1 NAND2X1_212 ( .A(wSelec[37]), .B(_1820_), .Y(_1827_) );
	NOR2X1 NOR2X1_117 ( .A(_1827_), .B(_1813_), .Y(_1828_) );
	NAND2X1 NAND2X1_213 ( .A(wData[32]), .B(_1828_), .Y(_1829_) );
	NAND2X1 NAND2X1_214 ( .A(wSelec[36]), .B(wSelec[37]), .Y(_1830_) );
	NOR2X1 NOR2X1_118 ( .A(_1830_), .B(_1817_), .Y(_1831_) );
	NOR2X1 NOR2X1_119 ( .A(_1830_), .B(_1808_), .Y(_1832_) );
	AOI22X1 AOI22X1_139 ( .A(_1831_), .B(wData[56]), .C(wData[52]), .D(_1832_), .Y(_1833_) );
	NOR2X1 NOR2X1_120 ( .A(_1823_), .B(_1830_), .Y(_1834_) );
	NOR2X1 NOR2X1_121 ( .A(_1823_), .B(_1827_), .Y(_1835_) );
	AOI22X1 AOI22X1_140 ( .A(wData[60]), .B(_1834_), .C(_1835_), .D(wData[44]), .Y(_1836_) );
	NAND3X1 NAND3X1_43 ( .A(_1829_), .B(_1836_), .C(_1833_), .Y(_1837_) );
	NOR2X1 NOR2X1_122 ( .A(_1817_), .B(_1827_), .Y(_1838_) );
	NAND2X1 NAND2X1_215 ( .A(wData[40]), .B(_1838_), .Y(_1839_) );
	NOR2X1 NOR2X1_123 ( .A(_1827_), .B(_1808_), .Y(_1840_) );
	NAND2X1 NAND2X1_216 ( .A(wData[36]), .B(_1840_), .Y(_1841_) );
	NOR2X1 NOR2X1_124 ( .A(_1821_), .B(_1813_), .Y(_1842_) );
	NAND2X1 NAND2X1_217 ( .A(wData[0]), .B(_1842_), .Y(_1843_) );
	NAND3X1 NAND3X1_44 ( .A(_1839_), .B(_1841_), .C(_1843_), .Y(_1844_) );
	INVX1 INVX1_125 ( .A(wData[48]), .Y(_1845_) );
	NOR2X1 NOR2X1_125 ( .A(_1820_), .B(_1809_), .Y(_1846_) );
	NAND2X1 NAND2X1_218 ( .A(_1812_), .B(_1846_), .Y(_1847_) );
	NOR2X1 NOR2X1_126 ( .A(_1817_), .B(_1821_), .Y(_1848_) );
	NOR2X1 NOR2X1_127 ( .A(_1823_), .B(_1821_), .Y(_1849_) );
	AOI22X1 AOI22X1_141 ( .A(_1848_), .B(wData[8]), .C(wData[12]), .D(_1849_), .Y(_1850_) );
	OAI21X1 OAI21X1_32 ( .A(_1845_), .B(_1847_), .C(_1850_), .Y(_1851_) );
	OR2X2 OR2X2_14 ( .A(_1851_), .B(_1844_), .Y(_1852_) );
	NOR3X1 NOR3X1_98 ( .A(_1826_), .B(_1837_), .C(_1852_), .Y(_1853_) );
	AND2X2 AND2X2_18 ( .A(_1853_), .B(_1617_), .Y(_1854_) );
	AOI21X1 AOI21X1_21 ( .A(_1708_), .B(_1806_), .C(_1854_), .Y(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_0_) );
	INVX1 INVX1_126 ( .A(_1725_), .Y(_1855_) );
	AOI21X1 AOI21X1_22 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_1855_), .C(_1617_), .Y(_1856_) );
	AOI22X1 AOI22X1_142 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_1625_), .C(_1641_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_1857_) );
	AOI22X1 AOI22X1_143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_1645_), .C(_1651_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_1858_) );
	NAND3X1 NAND3X1_45 ( .A(_1856_), .B(_1857_), .C(_1858_), .Y(_1859_) );
	INVX1 INVX1_127 ( .A(_1685_), .Y(_1860_) );
	AOI22X1 AOI22X1_144 ( .A(_1710_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_1860_), .Y(_1861_) );
	AOI22X1 AOI22X1_145 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_1784_), .C(_1663_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_1862_) );
	INVX1 INVX1_128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_1863_) );
	INVX1 INVX1_129 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_1864_) );
	OAI22X1 OAI22X1_26 ( .A(_1863_), .B(_1672_), .C(_1670_), .D(_1864_), .Y(_1865_) );
	INVX1 INVX1_130 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_1866_) );
	NAND2X1 NAND2X1_219 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_1773_), .Y(_1867_) );
	OAI21X1 OAI21X1_33 ( .A(_1866_), .B(_1678_), .C(_1867_), .Y(_1868_) );
	NOR2X1 NOR2X1_128 ( .A(_1865_), .B(_1868_), .Y(_1869_) );
	NAND3X1 NAND3X1_46 ( .A(_1861_), .B(_1862_), .C(_1869_), .Y(_1870_) );
	INVX1 INVX1_131 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_1871_) );
	NAND2X1 NAND2X1_220 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_1657_), .Y(_1872_) );
	OAI21X1 OAI21X1_34 ( .A(_1871_), .B(_1687_), .C(_1872_), .Y(_1873_) );
	INVX1 INVX1_132 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_1874_) );
	INVX1 INVX1_133 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_1875_) );
	OAI22X1 OAI22X1_27 ( .A(_1874_), .B(_1693_), .C(_1691_), .D(_1875_), .Y(_1876_) );
	NOR2X1 NOR2X1_129 ( .A(_1876_), .B(_1873_), .Y(_1877_) );
	AOI22X1 AOI22X1_146 ( .A(_1777_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_1750_), .Y(_1878_) );
	AND2X2 AND2X2_19 ( .A(_1624_), .B(_1639_), .Y(_1879_) );
	AOI22X1 AOI22X1_147 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_1749_), .C(_1879_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_1880_) );
	NAND3X1 NAND3X1_47 ( .A(_1878_), .B(_1880_), .C(_1877_), .Y(_1881_) );
	NOR3X1 NOR3X1_99 ( .A(_1881_), .B(_1859_), .C(_1870_), .Y(_1882_) );
	INVX1 INVX1_134 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_1883_) );
	NAND2X1 NAND2X1_221 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_1712_), .Y(_1884_) );
	OAI21X1 OAI21X1_35 ( .A(_1714_), .B(_1883_), .C(_1884_), .Y(_1885_) );
	AOI21X1 AOI21X1_23 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_1761_), .C(_1885_), .Y(_1886_) );
	INVX1 INVX1_135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_1887_) );
	INVX1 INVX1_136 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_1888_) );
	OAI22X1 OAI22X1_28 ( .A(_1888_), .B(_1720_), .C(_1721_), .D(_1887_), .Y(_1889_) );
	INVX1 INVX1_137 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_1890_) );
	NAND2X1 NAND2X1_222 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_1730_), .Y(_1891_) );
	OAI21X1 OAI21X1_36 ( .A(_1631_), .B(_1890_), .C(_1891_), .Y(_1892_) );
	NOR2X1 NOR2X1_130 ( .A(_1892_), .B(_1889_), .Y(_1893_) );
	INVX1 INVX1_138 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_1894_) );
	INVX1 INVX1_139 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_1895_) );
	OAI22X1 OAI22X1_29 ( .A(_1726_), .B(_1895_), .C(_1732_), .D(_1894_), .Y(_1896_) );
	INVX1 INVX1_140 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_1897_) );
	NOR2X1 NOR2X1_131 ( .A(_1897_), .B(_1737_), .Y(_1898_) );
	INVX1 INVX1_141 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_1899_) );
	NOR2X1 NOR2X1_132 ( .A(_1899_), .B(_1738_), .Y(_1900_) );
	NOR3X1 NOR3X1_100 ( .A(_1898_), .B(_1896_), .C(_1900_), .Y(_1901_) );
	NAND3X1 NAND3X1_48 ( .A(_1893_), .B(_1886_), .C(_1901_), .Y(_1902_) );
	AOI22X1 AOI22X1_148 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_1742_), .C(_1743_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_1903_) );
	AOI22X1 AOI22X1_149 ( .A(_1745_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_1746_), .Y(_1904_) );
	NAND2X1 NAND2X1_223 ( .A(_1903_), .B(_1904_), .Y(_1905_) );
	AOI22X1 AOI22X1_150 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_1753_), .C(_1752_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_1906_) );
	AOI22X1 AOI22X1_151 ( .A(_1696_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_1703_), .Y(_1907_) );
	NAND2X1 NAND2X1_224 ( .A(_1906_), .B(_1907_), .Y(_1908_) );
	NOR2X1 NOR2X1_133 ( .A(_1905_), .B(_1908_), .Y(_1909_) );
	AOI22X1 AOI22X1_152 ( .A(_1757_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_1758_), .Y(_1910_) );
	AOI22X1 AOI22X1_153 ( .A(_1659_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_1760_), .Y(_1911_) );
	NAND2X1 NAND2X1_225 ( .A(_1910_), .B(_1911_), .Y(_1912_) );
	AOI22X1 AOI22X1_154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_1764_), .C(_1765_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_1913_) );
	AOI22X1 AOI22X1_155 ( .A(_1767_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_1768_), .Y(_1914_) );
	NAND2X1 NAND2X1_226 ( .A(_1914_), .B(_1913_), .Y(_1915_) );
	NOR2X1 NOR2X1_134 ( .A(_1912_), .B(_1915_), .Y(_1916_) );
	NAND2X1 NAND2X1_227 ( .A(_1916_), .B(_1909_), .Y(_1917_) );
	AOI22X1 AOI22X1_156 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_1774_), .C(_1675_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_1918_) );
	AOI22X1 AOI22X1_157 ( .A(_1698_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_1776_), .Y(_1919_) );
	NAND2X1 NAND2X1_228 ( .A(_1918_), .B(_1919_), .Y(_1920_) );
	AOI22X1 AOI22X1_158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_1665_), .C(_1785_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_1921_) );
	NAND2X1 NAND2X1_229 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_1780_), .Y(_1922_) );
	NAND2X1 NAND2X1_230 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_1782_), .Y(_1923_) );
	NAND3X1 NAND3X1_49 ( .A(_1922_), .B(_1923_), .C(_1921_), .Y(_1924_) );
	NOR2X1 NOR2X1_135 ( .A(_1924_), .B(_1920_), .Y(_1925_) );
	AOI22X1 AOI22X1_159 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_1789_), .C(_1790_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_1926_) );
	NAND2X1 NAND2X1_231 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_1792_), .Y(_1927_) );
	NAND2X1 NAND2X1_232 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_1794_), .Y(_1928_) );
	NAND3X1 NAND3X1_50 ( .A(_1927_), .B(_1928_), .C(_1926_), .Y(_1929_) );
	AOI22X1 AOI22X1_160 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_1798_), .C(_1797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_1930_) );
	AOI22X1 AOI22X1_161 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_1801_), .C(_1800_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_1931_) );
	NAND2X1 NAND2X1_233 ( .A(_1930_), .B(_1931_), .Y(_1932_) );
	NOR2X1 NOR2X1_136 ( .A(_1932_), .B(_1929_), .Y(_1933_) );
	NAND2X1 NAND2X1_234 ( .A(_1925_), .B(_1933_), .Y(_1934_) );
	NOR3X1 NOR3X1_101 ( .A(_1917_), .B(_1902_), .C(_1934_), .Y(_1935_) );
	AOI21X1 AOI21X1_24 ( .A(wData[21]), .B(_1811_), .C(_1616_), .Y(_1936_) );
	AOI22X1 AOI22X1_162 ( .A(_1814_), .B(wData[17]), .C(wData[1]), .D(_1842_), .Y(_1937_) );
	AOI22X1 AOI22X1_163 ( .A(_1835_), .B(wData[45]), .C(wData[25]), .D(_1818_), .Y(_1938_) );
	NAND3X1 NAND3X1_51 ( .A(_1936_), .B(_1938_), .C(_1937_), .Y(_1939_) );
	NAND3X1 NAND3X1_52 ( .A(wData[49]), .B(_1812_), .C(_1846_), .Y(_1940_) );
	AOI22X1 AOI22X1_164 ( .A(wData[61]), .B(_1834_), .C(_1822_), .D(wData[5]), .Y(_1941_) );
	AND2X2 AND2X2_20 ( .A(_1941_), .B(_1940_), .Y(_1942_) );
	AOI22X1 AOI22X1_165 ( .A(_1831_), .B(wData[57]), .C(wData[41]), .D(_1838_), .Y(_1943_) );
	AOI22X1 AOI22X1_166 ( .A(wData[53]), .B(_1832_), .C(_1828_), .D(wData[33]), .Y(_1944_) );
	AND2X2 AND2X2_21 ( .A(_1944_), .B(_1943_), .Y(_1945_) );
	AOI22X1 AOI22X1_167 ( .A(_1848_), .B(wData[9]), .C(wData[13]), .D(_1849_), .Y(_1946_) );
	AOI22X1 AOI22X1_168 ( .A(_1824_), .B(wData[29]), .C(wData[37]), .D(_1840_), .Y(_1947_) );
	AND2X2 AND2X2_22 ( .A(_1946_), .B(_1947_), .Y(_1948_) );
	NAND3X1 NAND3X1_53 ( .A(_1942_), .B(_1948_), .C(_1945_), .Y(_1949_) );
	NOR2X1 NOR2X1_137 ( .A(_1939_), .B(_1949_), .Y(_1950_) );
	AOI21X1 AOI21X1_25 ( .A(_1882_), .B(_1935_), .C(_1950_), .Y(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_1_) );
	AOI21X1 AOI21X1_26 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_1855_), .C(_1617_), .Y(_1951_) );
	INVX1 INVX1_142 ( .A(_1714_), .Y(_1952_) );
	AOI22X1 AOI22X1_169 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_1625_), .C(_1952_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_1953_) );
	INVX1 INVX1_143 ( .A(_1726_), .Y(_1954_) );
	AOI22X1 AOI22X1_170 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_1761_), .C(_1954_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_1955_) );
	NAND3X1 NAND3X1_54 ( .A(_1955_), .B(_1951_), .C(_1953_), .Y(_1956_) );
	AOI22X1 AOI22X1_171 ( .A(_1710_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_1860_), .Y(_1957_) );
	AOI22X1 AOI22X1_172 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_1659_), .C(_1632_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_1958_) );
	INVX1 INVX1_144 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_1959_) );
	NAND2X1 NAND2X1_235 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_1749_), .Y(_1960_) );
	OAI21X1 OAI21X1_37 ( .A(_1959_), .B(_1721_), .C(_1960_), .Y(_1961_) );
	INVX1 INVX1_145 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_1962_) );
	NAND2X1 NAND2X1_236 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_1675_), .Y(_1963_) );
	OAI21X1 OAI21X1_38 ( .A(_1962_), .B(_1678_), .C(_1963_), .Y(_1964_) );
	NOR2X1 NOR2X1_138 ( .A(_1961_), .B(_1964_), .Y(_1965_) );
	NAND3X1 NAND3X1_55 ( .A(_1957_), .B(_1958_), .C(_1965_), .Y(_1966_) );
	INVX1 INVX1_146 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_1967_) );
	NAND2X1 NAND2X1_237 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_1657_), .Y(_1968_) );
	OAI21X1 OAI21X1_39 ( .A(_1967_), .B(_1687_), .C(_1968_), .Y(_1969_) );
	INVX1 INVX1_147 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_1970_) );
	INVX1 INVX1_148 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_1971_) );
	OAI22X1 OAI22X1_30 ( .A(_1970_), .B(_1693_), .C(_1691_), .D(_1971_), .Y(_1972_) );
	NOR2X1 NOR2X1_139 ( .A(_1972_), .B(_1969_), .Y(_1973_) );
	AOI22X1 AOI22X1_173 ( .A(_1777_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_1750_), .Y(_1974_) );
	AND2X2 AND2X2_23 ( .A(_1649_), .B(_1671_), .Y(_1975_) );
	AOI22X1 AOI22X1_174 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_1975_), .C(_1879_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_1976_) );
	NAND3X1 NAND3X1_56 ( .A(_1974_), .B(_1976_), .C(_1973_), .Y(_1977_) );
	NOR3X1 NOR3X1_102 ( .A(_1977_), .B(_1956_), .C(_1966_), .Y(_1978_) );
	INVX1 INVX1_149 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_1979_) );
	NOR3X1 NOR3X1_103 ( .A(_1979_), .B(_1644_), .C(_1643_), .Y(_1980_) );
	AND2X2 AND2X2_24 ( .A(_1665_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_1981_) );
	AND2X2 AND2X2_25 ( .A(_1785_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_1982_) );
	NOR3X1 NOR3X1_104 ( .A(_1982_), .B(_1981_), .C(_1980_), .Y(_1983_) );
	INVX1 INVX1_150 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_1984_) );
	INVX1 INVX1_151 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_1985_) );
	OAI22X1 OAI22X1_31 ( .A(_1985_), .B(_1720_), .C(_1670_), .D(_1984_), .Y(_1986_) );
	INVX1 INVX1_152 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_1987_) );
	INVX1 INVX1_153 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_1988_) );
	NAND2X1 NAND2X1_238 ( .A(_1661_), .B(_1662_), .Y(_1989_) );
	OAI22X1 OAI22X1_32 ( .A(_1989_), .B(_1988_), .C(_1987_), .D(_1640_), .Y(_1990_) );
	NOR2X1 NOR2X1_140 ( .A(_1986_), .B(_1990_), .Y(_1991_) );
	INVX1 INVX1_154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_1992_) );
	NOR3X1 NOR3X1_105 ( .A(_1621_), .B(_1638_), .C(_1629_), .Y(_1993_) );
	NAND2X1 NAND2X1_239 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_1993_), .Y(_1994_) );
	OAI21X1 OAI21X1_40 ( .A(_1650_), .B(_1992_), .C(_1994_), .Y(_1995_) );
	INVX1 INVX1_155 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_1996_) );
	INVX1 INVX1_156 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_1997_) );
	OAI22X1 OAI22X1_33 ( .A(_1737_), .B(_1997_), .C(_1996_), .D(_1738_), .Y(_1998_) );
	NOR2X1 NOR2X1_141 ( .A(_1995_), .B(_1998_), .Y(_1999_) );
	NAND3X1 NAND3X1_57 ( .A(_1983_), .B(_1999_), .C(_1991_), .Y(_2000_) );
	AOI22X1 AOI22X1_175 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_1742_), .C(_1743_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_2001_) );
	AOI22X1 AOI22X1_176 ( .A(_1745_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_1746_), .Y(_2002_) );
	NAND2X1 NAND2X1_240 ( .A(_2001_), .B(_2002_), .Y(_2003_) );
	AOI22X1 AOI22X1_177 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_1753_), .C(_1752_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_2004_) );
	AOI22X1 AOI22X1_178 ( .A(_1696_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_1703_), .Y(_2005_) );
	NAND2X1 NAND2X1_241 ( .A(_2004_), .B(_2005_), .Y(_2006_) );
	NOR2X1 NOR2X1_142 ( .A(_2003_), .B(_2006_), .Y(_2007_) );
	AOI22X1 AOI22X1_179 ( .A(_1757_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_1758_), .Y(_2008_) );
	AOI22X1 AOI22X1_180 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_1784_), .C(_1760_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_2009_) );
	NAND2X1 NAND2X1_242 ( .A(_2009_), .B(_2008_), .Y(_2010_) );
	AOI22X1 AOI22X1_181 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_1764_), .C(_1765_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_2011_) );
	AOI22X1 AOI22X1_182 ( .A(_1767_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_1768_), .Y(_2012_) );
	NAND2X1 NAND2X1_243 ( .A(_2012_), .B(_2011_), .Y(_2013_) );
	NOR2X1 NOR2X1_143 ( .A(_2010_), .B(_2013_), .Y(_2014_) );
	NAND2X1 NAND2X1_244 ( .A(_2014_), .B(_2007_), .Y(_2015_) );
	AOI22X1 AOI22X1_183 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_1774_), .C(_1773_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_2016_) );
	AOI22X1 AOI22X1_184 ( .A(_1698_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_1776_), .Y(_2017_) );
	NAND2X1 NAND2X1_245 ( .A(_2016_), .B(_2017_), .Y(_2018_) );
	AOI22X1 AOI22X1_185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_1782_), .C(_1780_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_2019_) );
	AOI22X1 AOI22X1_186 ( .A(_1712_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_1730_), .Y(_2020_) );
	NAND2X1 NAND2X1_246 ( .A(_2020_), .B(_2019_), .Y(_2021_) );
	NOR2X1 NOR2X1_144 ( .A(_2021_), .B(_2018_), .Y(_2022_) );
	AOI22X1 AOI22X1_187 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_1789_), .C(_1790_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_2023_) );
	NAND2X1 NAND2X1_247 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_1792_), .Y(_2024_) );
	NAND2X1 NAND2X1_248 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_1794_), .Y(_2025_) );
	NAND3X1 NAND3X1_58 ( .A(_2024_), .B(_2025_), .C(_2023_), .Y(_2026_) );
	AOI22X1 AOI22X1_188 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_1798_), .C(_1797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_2027_) );
	AOI22X1 AOI22X1_189 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_1801_), .C(_1800_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_2028_) );
	NAND2X1 NAND2X1_249 ( .A(_2027_), .B(_2028_), .Y(_2029_) );
	NOR2X1 NOR2X1_145 ( .A(_2029_), .B(_2026_), .Y(_2030_) );
	NAND2X1 NAND2X1_250 ( .A(_2022_), .B(_2030_), .Y(_2031_) );
	NOR3X1 NOR3X1_106 ( .A(_2015_), .B(_2000_), .C(_2031_), .Y(_2032_) );
	AOI22X1 AOI22X1_190 ( .A(_1838_), .B(wData[42]), .C(wData[38]), .D(_1840_), .Y(_2033_) );
	AOI22X1 AOI22X1_191 ( .A(_1835_), .B(wData[46]), .C(_1842_), .D(wData[2]), .Y(_2034_) );
	NAND2X1 NAND2X1_251 ( .A(_2033_), .B(_2034_), .Y(_2035_) );
	AOI21X1 AOI21X1_27 ( .A(wData[34]), .B(_1828_), .C(_2035_), .Y(_2036_) );
	INVX1 INVX1_157 ( .A(wData[50]), .Y(_2037_) );
	AOI22X1 AOI22X1_192 ( .A(_1848_), .B(wData[10]), .C(wData[14]), .D(_1849_), .Y(_2038_) );
	OAI21X1 OAI21X1_41 ( .A(_2037_), .B(_1847_), .C(_2038_), .Y(_2039_) );
	AOI22X1 AOI22X1_193 ( .A(_1811_), .B(wData[22]), .C(wData[18]), .D(_1814_), .Y(_2040_) );
	NAND2X1 NAND2X1_252 ( .A(wData[26]), .B(_1818_), .Y(_2041_) );
	AOI22X1 AOI22X1_194 ( .A(_1824_), .B(wData[30]), .C(wData[6]), .D(_1822_), .Y(_2042_) );
	NAND3X1 NAND3X1_59 ( .A(_2041_), .B(_2042_), .C(_2040_), .Y(_2043_) );
	NOR2X1 NOR2X1_146 ( .A(_2039_), .B(_2043_), .Y(_2044_) );
	NAND2X1 NAND2X1_253 ( .A(wData[58]), .B(_1831_), .Y(_2045_) );
	NAND2X1 NAND2X1_254 ( .A(wData[54]), .B(_1832_), .Y(_2046_) );
	NAND2X1 NAND2X1_255 ( .A(_2045_), .B(_2046_), .Y(_2047_) );
	AOI21X1 AOI21X1_28 ( .A(wData[62]), .B(_1834_), .C(_2047_), .Y(_2048_) );
	NAND3X1 NAND3X1_60 ( .A(_2036_), .B(_2048_), .C(_2044_), .Y(_2049_) );
	NOR2X1 NOR2X1_147 ( .A(_1616_), .B(_2049_), .Y(_2050_) );
	AOI21X1 AOI21X1_29 ( .A(_1978_), .B(_2032_), .C(_2050_), .Y(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_2_) );
	AOI21X1 AOI21X1_30 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_1860_), .C(_1617_), .Y(_2051_) );
	AOI22X1 AOI22X1_195 ( .A(_1632_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_1952_), .Y(_2052_) );
	AOI22X1 AOI22X1_196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_1954_), .C(_1710_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_2053_) );
	NAND3X1 NAND3X1_61 ( .A(_2053_), .B(_2051_), .C(_2052_), .Y(_2054_) );
	AOI22X1 AOI22X1_197 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_1659_), .C(_1657_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_2055_) );
	AOI22X1 AOI22X1_198 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_1730_), .C(_1855_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_2056_) );
	INVX1 INVX1_158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_2057_) );
	INVX1 INVX1_159 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_2058_) );
	OAI22X1 OAI22X1_34 ( .A(_2057_), .B(_1672_), .C(_1721_), .D(_2058_), .Y(_2059_) );
	INVX1 INVX1_160 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_2060_) );
	NAND2X1 NAND2X1_256 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_1773_), .Y(_2061_) );
	OAI21X1 OAI21X1_42 ( .A(_2060_), .B(_1678_), .C(_2061_), .Y(_2062_) );
	NOR2X1 NOR2X1_148 ( .A(_2059_), .B(_2062_), .Y(_2063_) );
	NAND3X1 NAND3X1_62 ( .A(_2055_), .B(_2056_), .C(_2063_), .Y(_2064_) );
	AND2X2 AND2X2_26 ( .A(_1686_), .B(_1620_), .Y(_2065_) );
	AOI22X1 AOI22X1_199 ( .A(_1625_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_2065_), .Y(_2066_) );
	AND2X2 AND2X2_27 ( .A(_1684_), .B(_1649_), .Y(_2067_) );
	AND2X2 AND2X2_28 ( .A(_1692_), .B(_1649_), .Y(_2068_) );
	AOI22X1 AOI22X1_200 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_2068_), .C(_2067_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_2069_) );
	NAND2X1 NAND2X1_257 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_1777_), .Y(_2070_) );
	NAND2X1 NAND2X1_258 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_1750_), .Y(_2071_) );
	NAND2X1 NAND2X1_259 ( .A(_2070_), .B(_2071_), .Y(_2072_) );
	INVX1 INVX1_161 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_2073_) );
	NAND2X1 NAND2X1_260 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_1749_), .Y(_2074_) );
	OAI21X1 OAI21X1_43 ( .A(_2073_), .B(_1702_), .C(_2074_), .Y(_2075_) );
	NOR2X1 NOR2X1_149 ( .A(_2072_), .B(_2075_), .Y(_2076_) );
	NAND3X1 NAND3X1_63 ( .A(_2066_), .B(_2069_), .C(_2076_), .Y(_2077_) );
	NOR3X1 NOR3X1_107 ( .A(_2064_), .B(_2054_), .C(_2077_), .Y(_2078_) );
	INVX1 INVX1_162 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_2079_) );
	NAND2X1 NAND2X1_261 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_1665_), .Y(_2080_) );
	OAI21X1 OAI21X1_44 ( .A(_1670_), .B(_2079_), .C(_2080_), .Y(_2081_) );
	AOI21X1 AOI21X1_31 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_1645_), .C(_2081_), .Y(_2082_) );
	INVX1 INVX1_163 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_2083_) );
	INVX1 INVX1_164 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_2084_) );
	OAI22X1 OAI22X1_35 ( .A(_1989_), .B(_2084_), .C(_2083_), .D(_1640_), .Y(_2085_) );
	INVX1 INVX1_165 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_2086_) );
	NAND2X1 NAND2X1_262 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_1785_), .Y(_2087_) );
	OAI21X1 OAI21X1_45 ( .A(_1650_), .B(_2086_), .C(_2087_), .Y(_2088_) );
	NOR2X1 NOR2X1_150 ( .A(_2088_), .B(_2085_), .Y(_2089_) );
	INVX1 INVX1_166 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_2090_) );
	INVX1 INVX1_167 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_2091_) );
	OAI22X1 OAI22X1_36 ( .A(_1737_), .B(_2091_), .C(_2090_), .D(_1738_), .Y(_2092_) );
	INVX1 INVX1_168 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_2093_) );
	NAND2X1 NAND2X1_263 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_1784_), .Y(_2094_) );
	OAI21X1 OAI21X1_46 ( .A(_2093_), .B(_1720_), .C(_2094_), .Y(_2095_) );
	NOR2X1 NOR2X1_151 ( .A(_2095_), .B(_2092_), .Y(_2096_) );
	NAND3X1 NAND3X1_64 ( .A(_2082_), .B(_2096_), .C(_2089_), .Y(_2097_) );
	AOI22X1 AOI22X1_201 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_1742_), .C(_1743_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_2098_) );
	AOI22X1 AOI22X1_202 ( .A(_1745_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_1746_), .Y(_2099_) );
	NAND2X1 NAND2X1_264 ( .A(_2098_), .B(_2099_), .Y(_2100_) );
	AOI22X1 AOI22X1_203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_1753_), .C(_1752_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_2101_) );
	AOI22X1 AOI22X1_204 ( .A(_1696_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_1703_), .Y(_2102_) );
	NAND2X1 NAND2X1_265 ( .A(_2101_), .B(_2102_), .Y(_2103_) );
	NOR2X1 NOR2X1_152 ( .A(_2100_), .B(_2103_), .Y(_2104_) );
	AOI22X1 AOI22X1_205 ( .A(_1757_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_1758_), .Y(_2105_) );
	AOI22X1 AOI22X1_206 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_1993_), .C(_1760_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_2106_) );
	NAND2X1 NAND2X1_266 ( .A(_2106_), .B(_2105_), .Y(_2107_) );
	AOI22X1 AOI22X1_207 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_1764_), .C(_1765_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_2108_) );
	AOI22X1 AOI22X1_208 ( .A(_1767_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_1768_), .Y(_2109_) );
	NAND2X1 NAND2X1_267 ( .A(_2109_), .B(_2108_), .Y(_2110_) );
	NOR2X1 NOR2X1_153 ( .A(_2107_), .B(_2110_), .Y(_2111_) );
	NAND2X1 NAND2X1_268 ( .A(_2111_), .B(_2104_), .Y(_2112_) );
	AOI22X1 AOI22X1_209 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_1774_), .C(_1675_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_2113_) );
	AOI22X1 AOI22X1_210 ( .A(_1698_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_1776_), .Y(_2114_) );
	NAND2X1 NAND2X1_269 ( .A(_2113_), .B(_2114_), .Y(_2115_) );
	AOI22X1 AOI22X1_211 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_1782_), .C(_1780_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_2116_) );
	AOI22X1 AOI22X1_212 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_1712_), .C(_1761_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_2117_) );
	NAND2X1 NAND2X1_270 ( .A(_2117_), .B(_2116_), .Y(_2118_) );
	NOR2X1 NOR2X1_154 ( .A(_2118_), .B(_2115_), .Y(_2119_) );
	AOI22X1 AOI22X1_213 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_1789_), .C(_1790_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_2120_) );
	NAND2X1 NAND2X1_271 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_1792_), .Y(_2121_) );
	NAND2X1 NAND2X1_272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_1794_), .Y(_2122_) );
	NAND3X1 NAND3X1_65 ( .A(_2121_), .B(_2122_), .C(_2120_), .Y(_2123_) );
	AOI22X1 AOI22X1_214 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_1798_), .C(_1797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_2124_) );
	AOI22X1 AOI22X1_215 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_1801_), .C(_1800_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_2125_) );
	NAND2X1 NAND2X1_273 ( .A(_2124_), .B(_2125_), .Y(_2126_) );
	NOR2X1 NOR2X1_155 ( .A(_2126_), .B(_2123_), .Y(_2127_) );
	NAND2X1 NAND2X1_274 ( .A(_2119_), .B(_2127_), .Y(_2128_) );
	NOR3X1 NOR3X1_108 ( .A(_2112_), .B(_2097_), .C(_2128_), .Y(_2129_) );
	NAND2X1 NAND2X1_275 ( .A(wData[59]), .B(_1831_), .Y(_2130_) );
	OAI21X1 OAI21X1_47 ( .A(_1615_), .B(wBusy_bF_buf0), .C(_2130_), .Y(_2131_) );
	NAND2X1 NAND2X1_276 ( .A(wData[7]), .B(_1822_), .Y(_2132_) );
	NAND2X1 NAND2X1_277 ( .A(wData[55]), .B(_1832_), .Y(_2133_) );
	AOI22X1 AOI22X1_216 ( .A(wData[63]), .B(_1834_), .C(_1824_), .D(wData[31]), .Y(_2134_) );
	NAND3X1 NAND3X1_66 ( .A(_2132_), .B(_2133_), .C(_2134_), .Y(_2135_) );
	OR2X2 OR2X2_15 ( .A(_2135_), .B(_2131_), .Y(_2136_) );
	INVX1 INVX1_169 ( .A(wData[51]), .Y(_2137_) );
	NAND2X1 NAND2X1_278 ( .A(wData[47]), .B(_1835_), .Y(_2138_) );
	OAI21X1 OAI21X1_48 ( .A(_2137_), .B(_1847_), .C(_2138_), .Y(_2139_) );
	AOI21X1 AOI21X1_32 ( .A(wData[3]), .B(_1842_), .C(_2139_), .Y(_2140_) );
	AOI22X1 AOI22X1_217 ( .A(_1848_), .B(wData[11]), .C(wData[15]), .D(_1849_), .Y(_2141_) );
	AOI22X1 AOI22X1_218 ( .A(_1811_), .B(wData[23]), .C(wData[27]), .D(_1818_), .Y(_2142_) );
	AND2X2 AND2X2_29 ( .A(_2141_), .B(_2142_), .Y(_2143_) );
	NAND2X1 NAND2X1_279 ( .A(wData[39]), .B(_1840_), .Y(_2144_) );
	NAND2X1 NAND2X1_280 ( .A(wData[43]), .B(_1838_), .Y(_2145_) );
	NAND2X1 NAND2X1_281 ( .A(_2144_), .B(_2145_), .Y(_2146_) );
	NAND2X1 NAND2X1_282 ( .A(wData[19]), .B(_1814_), .Y(_2147_) );
	NAND2X1 NAND2X1_283 ( .A(wData[35]), .B(_1828_), .Y(_2148_) );
	NAND2X1 NAND2X1_284 ( .A(_2147_), .B(_2148_), .Y(_2149_) );
	NOR2X1 NOR2X1_156 ( .A(_2146_), .B(_2149_), .Y(_2150_) );
	NAND3X1 NAND3X1_67 ( .A(_2143_), .B(_2140_), .C(_2150_), .Y(_2151_) );
	NOR2X1 NOR2X1_157 ( .A(_2136_), .B(_2151_), .Y(_2152_) );
	AOI21X1 AOI21X1_33 ( .A(_2078_), .B(_2129_), .C(_2152_), .Y(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_3_) );
	INVX1 INVX1_170 ( .A(wSelec[44]), .Y(_2153_) );
	NOR2X1 NOR2X1_158 ( .A(wBusy_bF_buf4), .B(_2153_), .Y(_2154_) );
	INVX1 INVX1_171 ( .A(_2154_), .Y(_2155_) );
	INVX1 INVX1_172 ( .A(wSelec[54]), .Y(_2156_) );
	NAND2X1 NAND2X1_285 ( .A(wSelec[53]), .B(_2156_), .Y(_2157_) );
	INVX2 INVX2_5 ( .A(_2157_), .Y(_2158_) );
	OR2X2 OR2X2_16 ( .A(wSelec[50]), .B(wSelec[49]), .Y(_2159_) );
	INVX1 INVX1_173 ( .A(wSelec[52]), .Y(_2160_) );
	NAND2X1 NAND2X1_286 ( .A(wSelec[51]), .B(_2160_), .Y(_2161_) );
	NOR2X1 NOR2X1_159 ( .A(_2159_), .B(_2161_), .Y(_2162_) );
	AND2X2 AND2X2_30 ( .A(_2162_), .B(_2158_), .Y(_2163_) );
	AOI21X1 AOI21X1_34 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_2163_), .C(_2155_), .Y(_2164_) );
	INVX1 INVX1_174 ( .A(wSelec[50]), .Y(_2165_) );
	NAND2X1 NAND2X1_287 ( .A(wSelec[49]), .B(_2165_), .Y(_2166_) );
	OR2X2 OR2X2_17 ( .A(wSelec[51]), .B(wSelec[52]), .Y(_2167_) );
	NOR2X1 NOR2X1_160 ( .A(_2167_), .B(_2166_), .Y(_2168_) );
	NAND2X1 NAND2X1_288 ( .A(_2158_), .B(_2168_), .Y(_2169_) );
	INVX1 INVX1_175 ( .A(_2169_), .Y(_2170_) );
	INVX1 INVX1_176 ( .A(wSelec[49]), .Y(_2171_) );
	NAND2X1 NAND2X1_289 ( .A(wSelec[50]), .B(_2171_), .Y(_2172_) );
	INVX1 INVX1_177 ( .A(wSelec[51]), .Y(_2173_) );
	NAND2X1 NAND2X1_290 ( .A(wSelec[52]), .B(_2173_), .Y(_2174_) );
	NOR2X1 NOR2X1_161 ( .A(_2172_), .B(_2174_), .Y(_2175_) );
	NAND2X1 NAND2X1_291 ( .A(wSelec[53]), .B(wSelec[54]), .Y(_2176_) );
	INVX1 INVX1_178 ( .A(_2176_), .Y(_2177_) );
	NAND2X1 NAND2X1_292 ( .A(_2177_), .B(_2175_), .Y(_2178_) );
	INVX1 INVX1_179 ( .A(_2178_), .Y(_2179_) );
	AOI22X1 AOI22X1_219 ( .A(_2170_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_2179_), .Y(_2180_) );
	OR2X2 OR2X2_18 ( .A(_2166_), .B(_2167_), .Y(_2181_) );
	OR2X2 OR2X2_19 ( .A(wSelec[53]), .B(wSelec[54]), .Y(_2182_) );
	NOR2X1 NOR2X1_162 ( .A(_2182_), .B(_2181_), .Y(_2183_) );
	NOR2X1 NOR2X1_163 ( .A(_2161_), .B(_2166_), .Y(_2184_) );
	INVX1 INVX1_180 ( .A(wSelec[53]), .Y(_2185_) );
	NAND2X1 NAND2X1_293 ( .A(wSelec[54]), .B(_2185_), .Y(_2186_) );
	INVX2 INVX2_6 ( .A(_2186_), .Y(_2187_) );
	NAND2X1 NAND2X1_294 ( .A(_2187_), .B(_2184_), .Y(_2188_) );
	INVX1 INVX1_181 ( .A(_2188_), .Y(_2189_) );
	AOI22X1 AOI22X1_220 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_2183_), .C(_2189_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_2190_) );
	NAND3X1 NAND3X1_68 ( .A(_2164_), .B(_2190_), .C(_2180_), .Y(_2191_) );
	NOR2X1 NOR2X1_164 ( .A(wSelec[50]), .B(wSelec[49]), .Y(_2192_) );
	NOR2X1 NOR2X1_165 ( .A(wSelec[51]), .B(wSelec[52]), .Y(_2193_) );
	NAND2X1 NAND2X1_295 ( .A(_2192_), .B(_2193_), .Y(_2194_) );
	NOR2X1 NOR2X1_166 ( .A(_2157_), .B(_2194_), .Y(_2195_) );
	NAND2X1 NAND2X1_296 ( .A(wSelec[50]), .B(wSelec[49]), .Y(_2196_) );
	NOR3X1 NOR3X1_109 ( .A(_2167_), .B(_2196_), .C(_2157_), .Y(_2197_) );
	AOI22X1 AOI22X1_221 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_2197_), .C(_2195_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_2198_) );
	INVX1 INVX1_182 ( .A(_2182_), .Y(_2199_) );
	NOR2X1 NOR2X1_167 ( .A(_2167_), .B(_2172_), .Y(_2200_) );
	AND2X2 AND2X2_31 ( .A(_2200_), .B(_2199_), .Y(_2201_) );
	NAND2X1 NAND2X1_297 ( .A(wSelec[51]), .B(wSelec[52]), .Y(_2202_) );
	NOR3X1 NOR3X1_110 ( .A(_2176_), .B(_2196_), .C(_2202_), .Y(_2203_) );
	AOI22X1 AOI22X1_222 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_2203_), .C(_2201_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_2204_) );
	INVX1 INVX1_183 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_2205_) );
	INVX1 INVX1_184 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_2206_) );
	NOR2X1 NOR2X1_168 ( .A(_2166_), .B(_2174_), .Y(_2207_) );
	NAND2X1 NAND2X1_298 ( .A(_2177_), .B(_2207_), .Y(_2208_) );
	NOR2X1 NOR2X1_169 ( .A(_2196_), .B(_2202_), .Y(_2209_) );
	NAND2X1 NAND2X1_299 ( .A(_2209_), .B(_2187_), .Y(_2210_) );
	OAI22X1 OAI22X1_37 ( .A(_2205_), .B(_2210_), .C(_2208_), .D(_2206_), .Y(_2211_) );
	INVX1 INVX1_185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_2212_) );
	NOR3X1 NOR3X1_111 ( .A(_2157_), .B(_2172_), .C(_2174_), .Y(_2213_) );
	NAND2X1 NAND2X1_300 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_2213_), .Y(_2214_) );
	NOR2X1 NOR2X1_170 ( .A(_2196_), .B(_2161_), .Y(_2215_) );
	NAND2X1 NAND2X1_301 ( .A(_2187_), .B(_2215_), .Y(_2216_) );
	OAI21X1 OAI21X1_49 ( .A(_2212_), .B(_2216_), .C(_2214_), .Y(_2217_) );
	NOR2X1 NOR2X1_171 ( .A(_2211_), .B(_2217_), .Y(_2218_) );
	NAND3X1 NAND3X1_69 ( .A(_2198_), .B(_2204_), .C(_2218_), .Y(_2219_) );
	INVX1 INVX1_186 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_2220_) );
	INVX1 INVX1_187 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_2221_) );
	NOR2X1 NOR2X1_172 ( .A(_2161_), .B(_2172_), .Y(_2222_) );
	NAND2X1 NAND2X1_302 ( .A(_2158_), .B(_2222_), .Y(_2223_) );
	NOR2X1 NOR2X1_173 ( .A(_2159_), .B(_2174_), .Y(_2224_) );
	NAND2X1 NAND2X1_303 ( .A(_2158_), .B(_2224_), .Y(_2225_) );
	OAI22X1 OAI22X1_38 ( .A(_2225_), .B(_2220_), .C(_2221_), .D(_2223_), .Y(_2226_) );
	INVX1 INVX1_188 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_2227_) );
	INVX1 INVX1_189 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_2228_) );
	NAND2X1 NAND2X1_304 ( .A(_2187_), .B(_2222_), .Y(_2229_) );
	NOR2X1 NOR2X1_174 ( .A(_2196_), .B(_2167_), .Y(_2230_) );
	NAND2X1 NAND2X1_305 ( .A(_2187_), .B(_2230_), .Y(_2231_) );
	OAI22X1 OAI22X1_39 ( .A(_2227_), .B(_2231_), .C(_2229_), .D(_2228_), .Y(_2232_) );
	NOR2X1 NOR2X1_175 ( .A(_2232_), .B(_2226_), .Y(_2233_) );
	NOR3X1 NOR3X1_112 ( .A(_2166_), .B(_2202_), .C(_2186_), .Y(_2234_) );
	NAND2X1 NAND2X1_306 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_2234_), .Y(_2235_) );
	NOR3X1 NOR3X1_113 ( .A(_2174_), .B(_2196_), .C(_2186_), .Y(_2236_) );
	NAND2X1 NAND2X1_307 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_2236_), .Y(_2237_) );
	NAND2X1 NAND2X1_308 ( .A(_2235_), .B(_2237_), .Y(_2238_) );
	INVX1 INVX1_190 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_2239_) );
	NAND2X1 NAND2X1_309 ( .A(_2177_), .B(_2162_), .Y(_2240_) );
	NOR3X1 NOR3X1_114 ( .A(_2172_), .B(_2174_), .C(_2186_), .Y(_2241_) );
	NAND2X1 NAND2X1_310 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_2241_), .Y(_2242_) );
	OAI21X1 OAI21X1_50 ( .A(_2239_), .B(_2240_), .C(_2242_), .Y(_2243_) );
	NOR2X1 NOR2X1_176 ( .A(_2238_), .B(_2243_), .Y(_2244_) );
	NAND2X1 NAND2X1_311 ( .A(_2233_), .B(_2244_), .Y(_2245_) );
	NOR3X1 NOR3X1_115 ( .A(_2191_), .B(_2245_), .C(_2219_), .Y(_2246_) );
	NAND2X1 NAND2X1_312 ( .A(_2158_), .B(_2215_), .Y(_2247_) );
	INVX1 INVX1_191 ( .A(_2247_), .Y(_2248_) );
	INVX1 INVX1_192 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_2249_) );
	NOR3X1 NOR3X1_116 ( .A(_2159_), .B(_2182_), .C(_2161_), .Y(_2250_) );
	NAND2X1 NAND2X1_313 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_2250_), .Y(_2251_) );
	NAND2X1 NAND2X1_314 ( .A(_2199_), .B(_2222_), .Y(_2252_) );
	OAI21X1 OAI21X1_51 ( .A(_2252_), .B(_2249_), .C(_2251_), .Y(_2253_) );
	AOI21X1 AOI21X1_35 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_2248_), .C(_2253_), .Y(_2254_) );
	INVX1 INVX1_193 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_2255_) );
	INVX1 INVX1_194 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_2256_) );
	NOR2X1 NOR2X1_177 ( .A(_2202_), .B(_2159_), .Y(_2257_) );
	NAND2X1 NAND2X1_315 ( .A(_2158_), .B(_2257_), .Y(_2258_) );
	NAND2X1 NAND2X1_316 ( .A(_2199_), .B(_2184_), .Y(_2259_) );
	OAI22X1 OAI22X1_40 ( .A(_2256_), .B(_2258_), .C(_2259_), .D(_2255_), .Y(_2260_) );
	INVX1 INVX1_195 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_2261_) );
	INVX1 INVX1_196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_2262_) );
	NAND2X1 NAND2X1_317 ( .A(_2158_), .B(_2184_), .Y(_2263_) );
	NAND2X1 NAND2X1_318 ( .A(_2199_), .B(_2230_), .Y(_2264_) );
	OAI22X1 OAI22X1_41 ( .A(_2261_), .B(_2264_), .C(_2263_), .D(_2262_), .Y(_2265_) );
	NOR2X1 NOR2X1_178 ( .A(_2260_), .B(_2265_), .Y(_2266_) );
	INVX1 INVX1_197 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_2267_) );
	NOR3X1 NOR3X1_117 ( .A(_2182_), .B(_2196_), .C(_2161_), .Y(_2268_) );
	NAND2X1 NAND2X1_319 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_2268_), .Y(_2269_) );
	OR2X2 OR2X2_20 ( .A(_2194_), .B(_2176_), .Y(_2270_) );
	OAI21X1 OAI21X1_52 ( .A(_2267_), .B(_2270_), .C(_2269_), .Y(_2271_) );
	INVX1 INVX1_198 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_2272_) );
	INVX1 INVX1_199 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_2273_) );
	NOR2X1 NOR2X1_179 ( .A(_2202_), .B(_2172_), .Y(_2274_) );
	NAND2X1 NAND2X1_320 ( .A(_2158_), .B(_2274_), .Y(_2275_) );
	NAND2X1 NAND2X1_321 ( .A(_2177_), .B(_2168_), .Y(_2276_) );
	OAI22X1 OAI22X1_42 ( .A(_2275_), .B(_2273_), .C(_2272_), .D(_2276_), .Y(_2277_) );
	NOR2X1 NOR2X1_180 ( .A(_2271_), .B(_2277_), .Y(_2278_) );
	NAND3X1 NAND3X1_70 ( .A(_2254_), .B(_2278_), .C(_2266_), .Y(_2279_) );
	NOR3X1 NOR3X1_118 ( .A(_2159_), .B(_2167_), .C(_2182_), .Y(_2280_) );
	NOR3X1 NOR3X1_119 ( .A(_2176_), .B(_2202_), .C(_2166_), .Y(_2281_) );
	AOI22X1 AOI22X1_223 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_2280_), .C(_2281_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_2282_) );
	NOR3X1 NOR3X1_120 ( .A(_2176_), .B(_2202_), .C(_2172_), .Y(_2283_) );
	NOR3X1 NOR3X1_121 ( .A(_2176_), .B(_2196_), .C(_2174_), .Y(_2284_) );
	AOI22X1 AOI22X1_224 ( .A(_2283_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_2284_), .Y(_2285_) );
	NAND2X1 NAND2X1_322 ( .A(_2282_), .B(_2285_), .Y(_2286_) );
	NOR3X1 NOR3X1_122 ( .A(_2174_), .B(_2159_), .C(_2186_), .Y(_2287_) );
	NOR3X1 NOR3X1_123 ( .A(_2166_), .B(_2174_), .C(_2186_), .Y(_2288_) );
	AOI22X1 AOI22X1_225 ( .A(_2287_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_2288_), .Y(_2289_) );
	NOR3X1 NOR3X1_124 ( .A(_2157_), .B(_2202_), .C(_2166_), .Y(_2290_) );
	NOR3X1 NOR3X1_125 ( .A(_2196_), .B(_2202_), .C(_2157_), .Y(_2291_) );
	AOI22X1 AOI22X1_226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_2291_), .C(_2290_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_2292_) );
	NAND2X1 NAND2X1_323 ( .A(_2292_), .B(_2289_), .Y(_2293_) );
	NOR2X1 NOR2X1_181 ( .A(_2286_), .B(_2293_), .Y(_2294_) );
	NOR3X1 NOR3X1_126 ( .A(_2182_), .B(_2202_), .C(_2166_), .Y(_2295_) );
	NOR3X1 NOR3X1_127 ( .A(_2182_), .B(_2202_), .C(_2172_), .Y(_2296_) );
	AOI22X1 AOI22X1_227 ( .A(_2295_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_2296_), .Y(_2297_) );
	NOR3X1 NOR3X1_128 ( .A(_2182_), .B(_2196_), .C(_2174_), .Y(_2298_) );
	NOR3X1 NOR3X1_129 ( .A(_2157_), .B(_2167_), .C(_2172_), .Y(_2299_) );
	AOI22X1 AOI22X1_228 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_2298_), .C(_2299_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_2300_) );
	NAND2X1 NAND2X1_324 ( .A(_2297_), .B(_2300_), .Y(_2301_) );
	NOR3X1 NOR3X1_130 ( .A(_2196_), .B(_2202_), .C(_2182_), .Y(_2302_) );
	NOR3X1 NOR3X1_131 ( .A(_2172_), .B(_2167_), .C(_2186_), .Y(_2303_) );
	AOI22X1 AOI22X1_229 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_2302_), .C(_2303_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_2304_) );
	NOR3X1 NOR3X1_132 ( .A(_2159_), .B(_2167_), .C(_2186_), .Y(_2305_) );
	NOR3X1 NOR3X1_133 ( .A(_2159_), .B(_2202_), .C(_2186_), .Y(_2306_) );
	AOI22X1 AOI22X1_230 ( .A(_2305_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_2306_), .Y(_2307_) );
	NAND2X1 NAND2X1_325 ( .A(_2307_), .B(_2304_), .Y(_2308_) );
	NOR2X1 NOR2X1_182 ( .A(_2301_), .B(_2308_), .Y(_2309_) );
	NAND2X1 NAND2X1_326 ( .A(_2309_), .B(_2294_), .Y(_2310_) );
	NOR3X1 NOR3X1_134 ( .A(_2157_), .B(_2196_), .C(_2174_), .Y(_2311_) );
	NOR3X1 NOR3X1_135 ( .A(_2167_), .B(_2176_), .C(_2172_), .Y(_2312_) );
	AOI22X1 AOI22X1_231 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_2312_), .C(_2311_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_2313_) );
	NOR3X1 NOR3X1_136 ( .A(_2161_), .B(_2159_), .C(_2186_), .Y(_2314_) );
	NOR3X1 NOR3X1_137 ( .A(_2172_), .B(_2202_), .C(_2186_), .Y(_2315_) );
	AOI22X1 AOI22X1_232 ( .A(_2314_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_2315_), .Y(_2316_) );
	NAND2X1 NAND2X1_327 ( .A(_2313_), .B(_2316_), .Y(_2317_) );
	NOR3X1 NOR3X1_138 ( .A(_2157_), .B(_2166_), .C(_2174_), .Y(_2318_) );
	NAND2X1 NAND2X1_328 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_2318_), .Y(_2319_) );
	NOR3X1 NOR3X1_139 ( .A(_2176_), .B(_2196_), .C(_2161_), .Y(_2320_) );
	NAND2X1 NAND2X1_329 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_2320_), .Y(_2321_) );
	NOR3X1 NOR3X1_140 ( .A(_2159_), .B(_2202_), .C(_2182_), .Y(_2322_) );
	NOR3X1 NOR3X1_141 ( .A(_2159_), .B(_2176_), .C(_2174_), .Y(_2323_) );
	AOI22X1 AOI22X1_233 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_2322_), .C(_2323_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_2324_) );
	NAND3X1 NAND3X1_71 ( .A(_2319_), .B(_2321_), .C(_2324_), .Y(_2325_) );
	NOR2X1 NOR2X1_183 ( .A(_2325_), .B(_2317_), .Y(_2326_) );
	NOR3X1 NOR3X1_142 ( .A(_2159_), .B(_2182_), .C(_2174_), .Y(_2327_) );
	NOR3X1 NOR3X1_143 ( .A(_2161_), .B(_2176_), .C(_2166_), .Y(_2328_) );
	AOI22X1 AOI22X1_234 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_2327_), .C(_2328_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_2329_) );
	NOR3X1 NOR3X1_144 ( .A(_2161_), .B(_2176_), .C(_2172_), .Y(_2330_) );
	NAND2X1 NAND2X1_330 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_2330_), .Y(_2331_) );
	NOR3X1 NOR3X1_145 ( .A(_2166_), .B(_2167_), .C(_2186_), .Y(_2332_) );
	NAND2X1 NAND2X1_331 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_2332_), .Y(_2333_) );
	NAND3X1 NAND3X1_72 ( .A(_2331_), .B(_2333_), .C(_2329_), .Y(_2334_) );
	NOR3X1 NOR3X1_146 ( .A(_2166_), .B(_2182_), .C(_2174_), .Y(_2335_) );
	NOR3X1 NOR3X1_147 ( .A(_2176_), .B(_2202_), .C(_2159_), .Y(_2336_) );
	AOI22X1 AOI22X1_235 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_2336_), .C(_2335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_2337_) );
	NOR3X1 NOR3X1_148 ( .A(_2172_), .B(_2182_), .C(_2174_), .Y(_2338_) );
	NOR3X1 NOR3X1_149 ( .A(_2176_), .B(_2196_), .C(_2167_), .Y(_2339_) );
	AOI22X1 AOI22X1_236 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_2339_), .C(_2338_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_2340_) );
	NAND2X1 NAND2X1_332 ( .A(_2337_), .B(_2340_), .Y(_2341_) );
	NOR2X1 NOR2X1_184 ( .A(_2341_), .B(_2334_), .Y(_2342_) );
	NAND2X1 NAND2X1_333 ( .A(_2326_), .B(_2342_), .Y(_2343_) );
	NOR3X1 NOR3X1_150 ( .A(_2310_), .B(_2279_), .C(_2343_), .Y(_2344_) );
	INVX1 INVX1_200 ( .A(wSelec[46]), .Y(_2345_) );
	NAND2X1 NAND2X1_334 ( .A(wSelec[45]), .B(_2345_), .Y(_2346_) );
	INVX1 INVX1_201 ( .A(wSelec[48]), .Y(_2347_) );
	NAND2X1 NAND2X1_335 ( .A(wSelec[47]), .B(_2347_), .Y(_2348_) );
	NOR2X1 NOR2X1_185 ( .A(_2346_), .B(_2348_), .Y(_2349_) );
	NOR2X1 NOR2X1_186 ( .A(wSelec[46]), .B(wSelec[45]), .Y(_2350_) );
	INVX1 INVX1_202 ( .A(_2350_), .Y(_2351_) );
	NOR2X1 NOR2X1_187 ( .A(_2348_), .B(_2351_), .Y(_2352_) );
	AOI22X1 AOI22X1_237 ( .A(wData[20]), .B(_2349_), .C(_2352_), .D(wData[16]), .Y(_2353_) );
	INVX1 INVX1_203 ( .A(wSelec[45]), .Y(_2354_) );
	NAND2X1 NAND2X1_336 ( .A(wSelec[46]), .B(_2354_), .Y(_2355_) );
	NOR2X1 NOR2X1_188 ( .A(_2355_), .B(_2348_), .Y(_2356_) );
	NAND2X1 NAND2X1_337 ( .A(wData[24]), .B(_2356_), .Y(_2357_) );
	INVX1 INVX1_204 ( .A(wSelec[47]), .Y(_2358_) );
	NAND2X1 NAND2X1_338 ( .A(_2358_), .B(_2347_), .Y(_2359_) );
	NOR2X1 NOR2X1_189 ( .A(_2346_), .B(_2359_), .Y(_2360_) );
	NAND2X1 NAND2X1_339 ( .A(wSelec[46]), .B(wSelec[45]), .Y(_2361_) );
	NOR2X1 NOR2X1_190 ( .A(_2361_), .B(_2348_), .Y(_2362_) );
	AOI22X1 AOI22X1_238 ( .A(_2362_), .B(wData[28]), .C(wData[4]), .D(_2360_), .Y(_2363_) );
	NAND3X1 NAND3X1_73 ( .A(_2357_), .B(_2363_), .C(_2353_), .Y(_2364_) );
	NAND2X1 NAND2X1_340 ( .A(wSelec[48]), .B(_2358_), .Y(_2365_) );
	NOR2X1 NOR2X1_191 ( .A(_2365_), .B(_2351_), .Y(_2366_) );
	NAND2X1 NAND2X1_341 ( .A(wData[32]), .B(_2366_), .Y(_2367_) );
	NAND2X1 NAND2X1_342 ( .A(wSelec[47]), .B(wSelec[48]), .Y(_2368_) );
	NOR2X1 NOR2X1_192 ( .A(_2368_), .B(_2355_), .Y(_2369_) );
	NOR2X1 NOR2X1_193 ( .A(_2368_), .B(_2346_), .Y(_2370_) );
	AOI22X1 AOI22X1_239 ( .A(_2369_), .B(wData[56]), .C(wData[52]), .D(_2370_), .Y(_2371_) );
	NOR2X1 NOR2X1_194 ( .A(_2361_), .B(_2368_), .Y(_2372_) );
	NOR2X1 NOR2X1_195 ( .A(_2361_), .B(_2365_), .Y(_2373_) );
	AOI22X1 AOI22X1_240 ( .A(wData[60]), .B(_2372_), .C(_2373_), .D(wData[44]), .Y(_2374_) );
	NAND3X1 NAND3X1_74 ( .A(_2367_), .B(_2374_), .C(_2371_), .Y(_2375_) );
	NOR2X1 NOR2X1_196 ( .A(_2355_), .B(_2365_), .Y(_2376_) );
	NAND2X1 NAND2X1_343 ( .A(wData[40]), .B(_2376_), .Y(_2377_) );
	NOR2X1 NOR2X1_197 ( .A(_2365_), .B(_2346_), .Y(_2378_) );
	NAND2X1 NAND2X1_344 ( .A(wData[36]), .B(_2378_), .Y(_2379_) );
	NOR2X1 NOR2X1_198 ( .A(_2359_), .B(_2351_), .Y(_2380_) );
	NAND2X1 NAND2X1_345 ( .A(wData[0]), .B(_2380_), .Y(_2381_) );
	NAND3X1 NAND3X1_75 ( .A(_2377_), .B(_2379_), .C(_2381_), .Y(_2382_) );
	INVX1 INVX1_205 ( .A(wData[48]), .Y(_2383_) );
	NOR2X1 NOR2X1_199 ( .A(_2358_), .B(_2347_), .Y(_2384_) );
	NAND2X1 NAND2X1_346 ( .A(_2350_), .B(_2384_), .Y(_2385_) );
	NOR2X1 NOR2X1_200 ( .A(_2355_), .B(_2359_), .Y(_2386_) );
	NOR2X1 NOR2X1_201 ( .A(_2361_), .B(_2359_), .Y(_2387_) );
	AOI22X1 AOI22X1_241 ( .A(_2386_), .B(wData[8]), .C(wData[12]), .D(_2387_), .Y(_2388_) );
	OAI21X1 OAI21X1_53 ( .A(_2383_), .B(_2385_), .C(_2388_), .Y(_2389_) );
	OR2X2 OR2X2_21 ( .A(_2389_), .B(_2382_), .Y(_2390_) );
	NOR3X1 NOR3X1_151 ( .A(_2364_), .B(_2375_), .C(_2390_), .Y(_2391_) );
	AND2X2 AND2X2_32 ( .A(_2391_), .B(_2155_), .Y(_2392_) );
	AOI21X1 AOI21X1_36 ( .A(_2246_), .B(_2344_), .C(_2392_), .Y(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_0_) );
	INVX1 INVX1_206 ( .A(_2263_), .Y(_2393_) );
	AOI21X1 AOI21X1_37 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_2393_), .C(_2155_), .Y(_2394_) );
	AOI22X1 AOI22X1_242 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_2163_), .C(_2179_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_2395_) );
	AOI22X1 AOI22X1_243 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_2183_), .C(_2189_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_2396_) );
	NAND3X1 NAND3X1_76 ( .A(_2394_), .B(_2395_), .C(_2396_), .Y(_2397_) );
	INVX1 INVX1_207 ( .A(_2223_), .Y(_2398_) );
	AOI22X1 AOI22X1_244 ( .A(_2248_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_2398_), .Y(_2399_) );
	AOI22X1 AOI22X1_245 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_2322_), .C(_2201_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_2400_) );
	INVX1 INVX1_208 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_2401_) );
	INVX1 INVX1_209 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_2402_) );
	OAI22X1 OAI22X1_43 ( .A(_2401_), .B(_2210_), .C(_2208_), .D(_2402_), .Y(_2403_) );
	INVX1 INVX1_210 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_2404_) );
	NAND2X1 NAND2X1_347 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_2311_), .Y(_2405_) );
	OAI21X1 OAI21X1_54 ( .A(_2404_), .B(_2216_), .C(_2405_), .Y(_2406_) );
	NOR2X1 NOR2X1_202 ( .A(_2403_), .B(_2406_), .Y(_2407_) );
	NAND3X1 NAND3X1_77 ( .A(_2399_), .B(_2400_), .C(_2407_), .Y(_2408_) );
	INVX1 INVX1_211 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_2409_) );
	NAND2X1 NAND2X1_348 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_2195_), .Y(_2410_) );
	OAI21X1 OAI21X1_55 ( .A(_2409_), .B(_2225_), .C(_2410_), .Y(_2411_) );
	INVX1 INVX1_212 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_2412_) );
	INVX1 INVX1_213 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_2413_) );
	OAI22X1 OAI22X1_44 ( .A(_2412_), .B(_2231_), .C(_2229_), .D(_2413_), .Y(_2414_) );
	NOR2X1 NOR2X1_203 ( .A(_2414_), .B(_2411_), .Y(_2415_) );
	AOI22X1 AOI22X1_246 ( .A(_2315_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_2288_), .Y(_2416_) );
	AND2X2 AND2X2_33 ( .A(_2162_), .B(_2177_), .Y(_2417_) );
	AOI22X1 AOI22X1_247 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_2287_), .C(_2417_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_2418_) );
	NAND3X1 NAND3X1_78 ( .A(_2416_), .B(_2418_), .C(_2415_), .Y(_2419_) );
	NOR3X1 NOR3X1_152 ( .A(_2419_), .B(_2397_), .C(_2408_), .Y(_2420_) );
	INVX1 INVX1_214 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_2421_) );
	NAND2X1 NAND2X1_349 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_2250_), .Y(_2422_) );
	OAI21X1 OAI21X1_56 ( .A(_2252_), .B(_2421_), .C(_2422_), .Y(_2423_) );
	AOI21X1 AOI21X1_38 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_2299_), .C(_2423_), .Y(_2424_) );
	INVX1 INVX1_215 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_2425_) );
	INVX1 INVX1_216 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_2426_) );
	OAI22X1 OAI22X1_45 ( .A(_2426_), .B(_2258_), .C(_2259_), .D(_2425_), .Y(_2427_) );
	INVX1 INVX1_217 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_2428_) );
	NAND2X1 NAND2X1_350 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_2268_), .Y(_2429_) );
	OAI21X1 OAI21X1_57 ( .A(_2169_), .B(_2428_), .C(_2429_), .Y(_2430_) );
	NOR2X1 NOR2X1_204 ( .A(_2430_), .B(_2427_), .Y(_2431_) );
	INVX1 INVX1_218 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_2432_) );
	INVX1 INVX1_219 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_2433_) );
	OAI22X1 OAI22X1_46 ( .A(_2264_), .B(_2433_), .C(_2270_), .D(_2432_), .Y(_2434_) );
	INVX1 INVX1_220 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_2435_) );
	NOR2X1 NOR2X1_205 ( .A(_2435_), .B(_2275_), .Y(_2436_) );
	INVX1 INVX1_221 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_2437_) );
	NOR2X1 NOR2X1_206 ( .A(_2437_), .B(_2276_), .Y(_2438_) );
	NOR3X1 NOR3X1_153 ( .A(_2436_), .B(_2434_), .C(_2438_), .Y(_2439_) );
	NAND3X1 NAND3X1_79 ( .A(_2431_), .B(_2424_), .C(_2439_), .Y(_2440_) );
	AOI22X1 AOI22X1_248 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_2280_), .C(_2281_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_2441_) );
	AOI22X1 AOI22X1_249 ( .A(_2283_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_2284_), .Y(_2442_) );
	NAND2X1 NAND2X1_351 ( .A(_2441_), .B(_2442_), .Y(_2443_) );
	AOI22X1 AOI22X1_250 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_2291_), .C(_2290_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_2444_) );
	AOI22X1 AOI22X1_251 ( .A(_2234_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_2241_), .Y(_2445_) );
	NAND2X1 NAND2X1_352 ( .A(_2444_), .B(_2445_), .Y(_2446_) );
	NOR2X1 NOR2X1_207 ( .A(_2443_), .B(_2446_), .Y(_2447_) );
	AOI22X1 AOI22X1_252 ( .A(_2295_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_2296_), .Y(_2448_) );
	AOI22X1 AOI22X1_253 ( .A(_2197_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_2298_), .Y(_2449_) );
	NAND2X1 NAND2X1_353 ( .A(_2448_), .B(_2449_), .Y(_2450_) );
	AOI22X1 AOI22X1_254 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_2302_), .C(_2303_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_2451_) );
	AOI22X1 AOI22X1_255 ( .A(_2305_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_2306_), .Y(_2452_) );
	NAND2X1 NAND2X1_354 ( .A(_2452_), .B(_2451_), .Y(_2453_) );
	NOR2X1 NOR2X1_208 ( .A(_2450_), .B(_2453_), .Y(_2454_) );
	NAND2X1 NAND2X1_355 ( .A(_2454_), .B(_2447_), .Y(_2455_) );
	AOI22X1 AOI22X1_256 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_2312_), .C(_2213_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_2456_) );
	AOI22X1 AOI22X1_257 ( .A(_2236_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_2314_), .Y(_2457_) );
	NAND2X1 NAND2X1_356 ( .A(_2456_), .B(_2457_), .Y(_2458_) );
	AOI22X1 AOI22X1_258 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_2203_), .C(_2323_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_2459_) );
	NAND2X1 NAND2X1_357 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_2318_), .Y(_2460_) );
	NAND2X1 NAND2X1_358 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_2320_), .Y(_2461_) );
	NAND3X1 NAND3X1_80 ( .A(_2460_), .B(_2461_), .C(_2459_), .Y(_2462_) );
	NOR2X1 NOR2X1_209 ( .A(_2462_), .B(_2458_), .Y(_2463_) );
	AOI22X1 AOI22X1_259 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_2327_), .C(_2328_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_2464_) );
	NAND2X1 NAND2X1_359 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_2330_), .Y(_2465_) );
	NAND2X1 NAND2X1_360 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_2332_), .Y(_2466_) );
	NAND3X1 NAND3X1_81 ( .A(_2465_), .B(_2466_), .C(_2464_), .Y(_2467_) );
	AOI22X1 AOI22X1_260 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_2336_), .C(_2335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_2468_) );
	AOI22X1 AOI22X1_261 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_2339_), .C(_2338_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_2469_) );
	NAND2X1 NAND2X1_361 ( .A(_2468_), .B(_2469_), .Y(_2470_) );
	NOR2X1 NOR2X1_210 ( .A(_2470_), .B(_2467_), .Y(_2471_) );
	NAND2X1 NAND2X1_362 ( .A(_2463_), .B(_2471_), .Y(_2472_) );
	NOR3X1 NOR3X1_154 ( .A(_2455_), .B(_2440_), .C(_2472_), .Y(_2473_) );
	AOI21X1 AOI21X1_39 ( .A(wData[21]), .B(_2349_), .C(_2154_), .Y(_2474_) );
	AOI22X1 AOI22X1_262 ( .A(_2352_), .B(wData[17]), .C(wData[1]), .D(_2380_), .Y(_2475_) );
	AOI22X1 AOI22X1_263 ( .A(_2373_), .B(wData[45]), .C(wData[25]), .D(_2356_), .Y(_2476_) );
	NAND3X1 NAND3X1_82 ( .A(_2474_), .B(_2476_), .C(_2475_), .Y(_2477_) );
	NAND3X1 NAND3X1_83 ( .A(wData[49]), .B(_2350_), .C(_2384_), .Y(_2478_) );
	AOI22X1 AOI22X1_264 ( .A(wData[61]), .B(_2372_), .C(_2360_), .D(wData[5]), .Y(_2479_) );
	AND2X2 AND2X2_34 ( .A(_2479_), .B(_2478_), .Y(_2480_) );
	AOI22X1 AOI22X1_265 ( .A(_2369_), .B(wData[57]), .C(wData[41]), .D(_2376_), .Y(_2481_) );
	AOI22X1 AOI22X1_266 ( .A(wData[53]), .B(_2370_), .C(_2366_), .D(wData[33]), .Y(_2482_) );
	AND2X2 AND2X2_35 ( .A(_2482_), .B(_2481_), .Y(_2483_) );
	AOI22X1 AOI22X1_267 ( .A(_2386_), .B(wData[9]), .C(wData[13]), .D(_2387_), .Y(_2484_) );
	AOI22X1 AOI22X1_268 ( .A(_2362_), .B(wData[29]), .C(wData[37]), .D(_2378_), .Y(_2485_) );
	AND2X2 AND2X2_36 ( .A(_2484_), .B(_2485_), .Y(_2486_) );
	NAND3X1 NAND3X1_84 ( .A(_2480_), .B(_2486_), .C(_2483_), .Y(_2487_) );
	NOR2X1 NOR2X1_211 ( .A(_2477_), .B(_2487_), .Y(_2488_) );
	AOI21X1 AOI21X1_40 ( .A(_2420_), .B(_2473_), .C(_2488_), .Y(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_1_) );
	AOI21X1 AOI21X1_41 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_2393_), .C(_2155_), .Y(_2489_) );
	INVX1 INVX1_222 ( .A(_2252_), .Y(_2490_) );
	AOI22X1 AOI22X1_269 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_2163_), .C(_2490_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_2491_) );
	INVX1 INVX1_223 ( .A(_2264_), .Y(_2492_) );
	AOI22X1 AOI22X1_270 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_2299_), .C(_2492_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_2493_) );
	NAND3X1 NAND3X1_85 ( .A(_2493_), .B(_2489_), .C(_2491_), .Y(_2494_) );
	AOI22X1 AOI22X1_271 ( .A(_2248_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_2398_), .Y(_2495_) );
	AOI22X1 AOI22X1_272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_2197_), .C(_2170_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_2496_) );
	INVX1 INVX1_224 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_2497_) );
	NAND2X1 NAND2X1_363 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_2287_), .Y(_2498_) );
	OAI21X1 OAI21X1_58 ( .A(_2497_), .B(_2259_), .C(_2498_), .Y(_2499_) );
	INVX1 INVX1_225 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_2500_) );
	NAND2X1 NAND2X1_364 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_2213_), .Y(_2501_) );
	OAI21X1 OAI21X1_59 ( .A(_2500_), .B(_2216_), .C(_2501_), .Y(_2502_) );
	NOR2X1 NOR2X1_212 ( .A(_2499_), .B(_2502_), .Y(_2503_) );
	NAND3X1 NAND3X1_86 ( .A(_2495_), .B(_2496_), .C(_2503_), .Y(_2504_) );
	INVX1 INVX1_226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_2505_) );
	NAND2X1 NAND2X1_365 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_2195_), .Y(_2506_) );
	OAI21X1 OAI21X1_60 ( .A(_2505_), .B(_2225_), .C(_2506_), .Y(_2507_) );
	INVX1 INVX1_227 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_2508_) );
	INVX1 INVX1_228 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_2509_) );
	OAI22X1 OAI22X1_47 ( .A(_2508_), .B(_2231_), .C(_2229_), .D(_2509_), .Y(_2510_) );
	NOR2X1 NOR2X1_213 ( .A(_2510_), .B(_2507_), .Y(_2511_) );
	AOI22X1 AOI22X1_273 ( .A(_2315_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_2288_), .Y(_2512_) );
	AND2X2 AND2X2_37 ( .A(_2187_), .B(_2209_), .Y(_2513_) );
	AOI22X1 AOI22X1_274 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_2513_), .C(_2417_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_2514_) );
	NAND3X1 NAND3X1_87 ( .A(_2512_), .B(_2514_), .C(_2511_), .Y(_2515_) );
	NOR3X1 NOR3X1_155 ( .A(_2515_), .B(_2494_), .C(_2504_), .Y(_2516_) );
	INVX1 INVX1_229 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_2517_) );
	NOR3X1 NOR3X1_156 ( .A(_2517_), .B(_2182_), .C(_2181_), .Y(_2518_) );
	AND2X2 AND2X2_38 ( .A(_2203_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_2519_) );
	AND2X2 AND2X2_39 ( .A(_2323_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_2520_) );
	NOR3X1 NOR3X1_157 ( .A(_2520_), .B(_2519_), .C(_2518_), .Y(_2521_) );
	INVX1 INVX1_230 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_2522_) );
	INVX1 INVX1_231 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_2523_) );
	OAI22X1 OAI22X1_48 ( .A(_2523_), .B(_2258_), .C(_2208_), .D(_2522_), .Y(_2524_) );
	INVX1 INVX1_232 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_2525_) );
	INVX1 INVX1_233 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_2526_) );
	NAND2X1 NAND2X1_366 ( .A(_2199_), .B(_2200_), .Y(_2527_) );
	OAI22X1 OAI22X1_49 ( .A(_2527_), .B(_2526_), .C(_2525_), .D(_2178_), .Y(_2528_) );
	NOR2X1 NOR2X1_214 ( .A(_2524_), .B(_2528_), .Y(_2529_) );
	INVX1 INVX1_234 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_2530_) );
	NOR3X1 NOR3X1_158 ( .A(_2159_), .B(_2176_), .C(_2167_), .Y(_2531_) );
	NAND2X1 NAND2X1_367 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_2531_), .Y(_2532_) );
	OAI21X1 OAI21X1_61 ( .A(_2188_), .B(_2530_), .C(_2532_), .Y(_2533_) );
	INVX1 INVX1_235 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_2534_) );
	INVX1 INVX1_236 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_2535_) );
	OAI22X1 OAI22X1_50 ( .A(_2275_), .B(_2535_), .C(_2534_), .D(_2276_), .Y(_2536_) );
	NOR2X1 NOR2X1_215 ( .A(_2533_), .B(_2536_), .Y(_2537_) );
	NAND3X1 NAND3X1_88 ( .A(_2521_), .B(_2537_), .C(_2529_), .Y(_2538_) );
	AOI22X1 AOI22X1_275 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_2280_), .C(_2281_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_2539_) );
	AOI22X1 AOI22X1_276 ( .A(_2283_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_2284_), .Y(_2540_) );
	NAND2X1 NAND2X1_368 ( .A(_2539_), .B(_2540_), .Y(_2541_) );
	AOI22X1 AOI22X1_277 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_2291_), .C(_2290_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_2542_) );
	AOI22X1 AOI22X1_278 ( .A(_2234_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_2241_), .Y(_2543_) );
	NAND2X1 NAND2X1_369 ( .A(_2542_), .B(_2543_), .Y(_2544_) );
	NOR2X1 NOR2X1_216 ( .A(_2541_), .B(_2544_), .Y(_2545_) );
	AOI22X1 AOI22X1_279 ( .A(_2295_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_2296_), .Y(_2546_) );
	AOI22X1 AOI22X1_280 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_2322_), .C(_2298_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_2547_) );
	NAND2X1 NAND2X1_370 ( .A(_2547_), .B(_2546_), .Y(_2548_) );
	AOI22X1 AOI22X1_281 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_2302_), .C(_2303_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_2549_) );
	AOI22X1 AOI22X1_282 ( .A(_2305_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_2306_), .Y(_2550_) );
	NAND2X1 NAND2X1_371 ( .A(_2550_), .B(_2549_), .Y(_2551_) );
	NOR2X1 NOR2X1_217 ( .A(_2548_), .B(_2551_), .Y(_2552_) );
	NAND2X1 NAND2X1_372 ( .A(_2552_), .B(_2545_), .Y(_2553_) );
	AOI22X1 AOI22X1_283 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_2312_), .C(_2311_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_2554_) );
	AOI22X1 AOI22X1_284 ( .A(_2236_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_2314_), .Y(_2555_) );
	NAND2X1 NAND2X1_373 ( .A(_2554_), .B(_2555_), .Y(_2556_) );
	AOI22X1 AOI22X1_285 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_2320_), .C(_2318_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_2557_) );
	AOI22X1 AOI22X1_286 ( .A(_2250_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_2268_), .Y(_2558_) );
	NAND2X1 NAND2X1_374 ( .A(_2558_), .B(_2557_), .Y(_2559_) );
	NOR2X1 NOR2X1_218 ( .A(_2559_), .B(_2556_), .Y(_2560_) );
	AOI22X1 AOI22X1_287 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_2327_), .C(_2328_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_2561_) );
	NAND2X1 NAND2X1_375 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_2330_), .Y(_2562_) );
	NAND2X1 NAND2X1_376 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_2332_), .Y(_2563_) );
	NAND3X1 NAND3X1_89 ( .A(_2562_), .B(_2563_), .C(_2561_), .Y(_2564_) );
	AOI22X1 AOI22X1_288 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_2336_), .C(_2335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_2565_) );
	AOI22X1 AOI22X1_289 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_2339_), .C(_2338_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_2566_) );
	NAND2X1 NAND2X1_377 ( .A(_2565_), .B(_2566_), .Y(_2567_) );
	NOR2X1 NOR2X1_219 ( .A(_2567_), .B(_2564_), .Y(_2568_) );
	NAND2X1 NAND2X1_378 ( .A(_2560_), .B(_2568_), .Y(_2569_) );
	NOR3X1 NOR3X1_159 ( .A(_2553_), .B(_2538_), .C(_2569_), .Y(_2570_) );
	AOI22X1 AOI22X1_290 ( .A(_2376_), .B(wData[42]), .C(wData[38]), .D(_2378_), .Y(_2571_) );
	AOI22X1 AOI22X1_291 ( .A(_2373_), .B(wData[46]), .C(_2380_), .D(wData[2]), .Y(_2572_) );
	NAND2X1 NAND2X1_379 ( .A(_2571_), .B(_2572_), .Y(_2573_) );
	AOI21X1 AOI21X1_42 ( .A(wData[34]), .B(_2366_), .C(_2573_), .Y(_2574_) );
	INVX1 INVX1_237 ( .A(wData[50]), .Y(_2575_) );
	AOI22X1 AOI22X1_292 ( .A(_2386_), .B(wData[10]), .C(wData[14]), .D(_2387_), .Y(_2576_) );
	OAI21X1 OAI21X1_62 ( .A(_2575_), .B(_2385_), .C(_2576_), .Y(_2577_) );
	AOI22X1 AOI22X1_293 ( .A(_2349_), .B(wData[22]), .C(wData[18]), .D(_2352_), .Y(_2578_) );
	NAND2X1 NAND2X1_380 ( .A(wData[26]), .B(_2356_), .Y(_2579_) );
	AOI22X1 AOI22X1_294 ( .A(_2362_), .B(wData[30]), .C(wData[6]), .D(_2360_), .Y(_2580_) );
	NAND3X1 NAND3X1_90 ( .A(_2579_), .B(_2580_), .C(_2578_), .Y(_2581_) );
	NOR2X1 NOR2X1_220 ( .A(_2577_), .B(_2581_), .Y(_2582_) );
	NAND2X1 NAND2X1_381 ( .A(wData[58]), .B(_2369_), .Y(_2583_) );
	NAND2X1 NAND2X1_382 ( .A(wData[54]), .B(_2370_), .Y(_2584_) );
	NAND2X1 NAND2X1_383 ( .A(_2583_), .B(_2584_), .Y(_2585_) );
	AOI21X1 AOI21X1_43 ( .A(wData[62]), .B(_2372_), .C(_2585_), .Y(_2586_) );
	NAND3X1 NAND3X1_91 ( .A(_2574_), .B(_2586_), .C(_2582_), .Y(_2587_) );
	NOR2X1 NOR2X1_221 ( .A(_2154_), .B(_2587_), .Y(_2588_) );
	AOI21X1 AOI21X1_44 ( .A(_2516_), .B(_2570_), .C(_2588_), .Y(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_2_) );
	AOI21X1 AOI21X1_45 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_2398_), .C(_2155_), .Y(_2589_) );
	AOI22X1 AOI22X1_295 ( .A(_2170_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_2490_), .Y(_2590_) );
	AOI22X1 AOI22X1_296 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_2492_), .C(_2248_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_2591_) );
	NAND3X1 NAND3X1_92 ( .A(_2591_), .B(_2589_), .C(_2590_), .Y(_2592_) );
	AOI22X1 AOI22X1_297 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_2197_), .C(_2195_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_2593_) );
	AOI22X1 AOI22X1_298 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_2268_), .C(_2393_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_2594_) );
	INVX1 INVX1_238 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_2595_) );
	INVX1 INVX1_239 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_2596_) );
	OAI22X1 OAI22X1_51 ( .A(_2595_), .B(_2210_), .C(_2259_), .D(_2596_), .Y(_2597_) );
	INVX1 INVX1_240 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_2598_) );
	NAND2X1 NAND2X1_384 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_2311_), .Y(_2599_) );
	OAI21X1 OAI21X1_63 ( .A(_2598_), .B(_2216_), .C(_2599_), .Y(_2600_) );
	NOR2X1 NOR2X1_222 ( .A(_2597_), .B(_2600_), .Y(_2601_) );
	NAND3X1 NAND3X1_93 ( .A(_2593_), .B(_2594_), .C(_2601_), .Y(_2602_) );
	AND2X2 AND2X2_40 ( .A(_2224_), .B(_2158_), .Y(_2603_) );
	AOI22X1 AOI22X1_299 ( .A(_2163_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_2603_), .Y(_2604_) );
	AND2X2 AND2X2_41 ( .A(_2222_), .B(_2187_), .Y(_2605_) );
	AND2X2 AND2X2_42 ( .A(_2230_), .B(_2187_), .Y(_2606_) );
	AOI22X1 AOI22X1_300 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_2606_), .C(_2605_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_2607_) );
	NAND2X1 NAND2X1_385 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_2315_), .Y(_2608_) );
	NAND2X1 NAND2X1_386 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_2288_), .Y(_2609_) );
	NAND2X1 NAND2X1_387 ( .A(_2608_), .B(_2609_), .Y(_2610_) );
	INVX1 INVX1_241 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_2611_) );
	NAND2X1 NAND2X1_388 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_2287_), .Y(_2612_) );
	OAI21X1 OAI21X1_64 ( .A(_2611_), .B(_2240_), .C(_2612_), .Y(_2613_) );
	NOR2X1 NOR2X1_223 ( .A(_2610_), .B(_2613_), .Y(_2614_) );
	NAND3X1 NAND3X1_94 ( .A(_2604_), .B(_2607_), .C(_2614_), .Y(_2615_) );
	NOR3X1 NOR3X1_160 ( .A(_2602_), .B(_2592_), .C(_2615_), .Y(_2616_) );
	INVX1 INVX1_242 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_2617_) );
	NAND2X1 NAND2X1_389 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_2203_), .Y(_2618_) );
	OAI21X1 OAI21X1_65 ( .A(_2208_), .B(_2617_), .C(_2618_), .Y(_2619_) );
	AOI21X1 AOI21X1_46 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_2183_), .C(_2619_), .Y(_2620_) );
	INVX1 INVX1_243 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_2621_) );
	INVX1 INVX1_244 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_2622_) );
	OAI22X1 OAI22X1_52 ( .A(_2527_), .B(_2622_), .C(_2621_), .D(_2178_), .Y(_2623_) );
	INVX1 INVX1_245 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_2624_) );
	NAND2X1 NAND2X1_390 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_2323_), .Y(_2625_) );
	OAI21X1 OAI21X1_66 ( .A(_2188_), .B(_2624_), .C(_2625_), .Y(_2626_) );
	NOR2X1 NOR2X1_224 ( .A(_2626_), .B(_2623_), .Y(_2627_) );
	INVX1 INVX1_246 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_2628_) );
	INVX1 INVX1_247 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_2629_) );
	OAI22X1 OAI22X1_53 ( .A(_2275_), .B(_2629_), .C(_2628_), .D(_2276_), .Y(_2630_) );
	INVX1 INVX1_248 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_2631_) );
	NAND2X1 NAND2X1_391 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_2322_), .Y(_2632_) );
	OAI21X1 OAI21X1_67 ( .A(_2631_), .B(_2258_), .C(_2632_), .Y(_2633_) );
	NOR2X1 NOR2X1_225 ( .A(_2633_), .B(_2630_), .Y(_2634_) );
	NAND3X1 NAND3X1_95 ( .A(_2620_), .B(_2634_), .C(_2627_), .Y(_2635_) );
	AOI22X1 AOI22X1_301 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_2280_), .C(_2281_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_2636_) );
	AOI22X1 AOI22X1_302 ( .A(_2283_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_2284_), .Y(_2637_) );
	NAND2X1 NAND2X1_392 ( .A(_2636_), .B(_2637_), .Y(_2638_) );
	AOI22X1 AOI22X1_303 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_2291_), .C(_2290_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_2639_) );
	AOI22X1 AOI22X1_304 ( .A(_2234_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_2241_), .Y(_2640_) );
	NAND2X1 NAND2X1_393 ( .A(_2639_), .B(_2640_), .Y(_2641_) );
	NOR2X1 NOR2X1_226 ( .A(_2638_), .B(_2641_), .Y(_2642_) );
	AOI22X1 AOI22X1_305 ( .A(_2295_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_2296_), .Y(_2643_) );
	AOI22X1 AOI22X1_306 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_2531_), .C(_2298_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_2644_) );
	NAND2X1 NAND2X1_394 ( .A(_2644_), .B(_2643_), .Y(_2645_) );
	AOI22X1 AOI22X1_307 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_2302_), .C(_2303_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_2646_) );
	AOI22X1 AOI22X1_308 ( .A(_2305_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_2306_), .Y(_2647_) );
	NAND2X1 NAND2X1_395 ( .A(_2647_), .B(_2646_), .Y(_2648_) );
	NOR2X1 NOR2X1_227 ( .A(_2645_), .B(_2648_), .Y(_2649_) );
	NAND2X1 NAND2X1_396 ( .A(_2649_), .B(_2642_), .Y(_2650_) );
	AOI22X1 AOI22X1_309 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_2312_), .C(_2213_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_2651_) );
	AOI22X1 AOI22X1_310 ( .A(_2236_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_2314_), .Y(_2652_) );
	NAND2X1 NAND2X1_397 ( .A(_2651_), .B(_2652_), .Y(_2653_) );
	AOI22X1 AOI22X1_311 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_2320_), .C(_2318_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_2654_) );
	AOI22X1 AOI22X1_312 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_2250_), .C(_2299_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_2655_) );
	NAND2X1 NAND2X1_398 ( .A(_2655_), .B(_2654_), .Y(_2656_) );
	NOR2X1 NOR2X1_228 ( .A(_2656_), .B(_2653_), .Y(_2657_) );
	AOI22X1 AOI22X1_313 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_2327_), .C(_2328_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_2658_) );
	NAND2X1 NAND2X1_399 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_2330_), .Y(_2659_) );
	NAND2X1 NAND2X1_400 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_2332_), .Y(_2660_) );
	NAND3X1 NAND3X1_96 ( .A(_2659_), .B(_2660_), .C(_2658_), .Y(_2661_) );
	AOI22X1 AOI22X1_314 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_2336_), .C(_2335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_2662_) );
	AOI22X1 AOI22X1_315 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_2339_), .C(_2338_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_2663_) );
	NAND2X1 NAND2X1_401 ( .A(_2662_), .B(_2663_), .Y(_2664_) );
	NOR2X1 NOR2X1_229 ( .A(_2664_), .B(_2661_), .Y(_2665_) );
	NAND2X1 NAND2X1_402 ( .A(_2657_), .B(_2665_), .Y(_2666_) );
	NOR3X1 NOR3X1_161 ( .A(_2650_), .B(_2635_), .C(_2666_), .Y(_2667_) );
	NAND2X1 NAND2X1_403 ( .A(wData[59]), .B(_2369_), .Y(_2668_) );
	OAI21X1 OAI21X1_68 ( .A(_2153_), .B(wBusy_bF_buf3), .C(_2668_), .Y(_2669_) );
	NAND2X1 NAND2X1_404 ( .A(wData[7]), .B(_2360_), .Y(_2670_) );
	NAND2X1 NAND2X1_405 ( .A(wData[55]), .B(_2370_), .Y(_2671_) );
	AOI22X1 AOI22X1_316 ( .A(wData[63]), .B(_2372_), .C(_2362_), .D(wData[31]), .Y(_2672_) );
	NAND3X1 NAND3X1_97 ( .A(_2670_), .B(_2671_), .C(_2672_), .Y(_2673_) );
	OR2X2 OR2X2_22 ( .A(_2673_), .B(_2669_), .Y(_2674_) );
	INVX1 INVX1_249 ( .A(wData[51]), .Y(_2675_) );
	NAND2X1 NAND2X1_406 ( .A(wData[47]), .B(_2373_), .Y(_2676_) );
	OAI21X1 OAI21X1_69 ( .A(_2675_), .B(_2385_), .C(_2676_), .Y(_2677_) );
	AOI21X1 AOI21X1_47 ( .A(wData[3]), .B(_2380_), .C(_2677_), .Y(_2678_) );
	AOI22X1 AOI22X1_317 ( .A(_2386_), .B(wData[11]), .C(wData[15]), .D(_2387_), .Y(_2679_) );
	AOI22X1 AOI22X1_318 ( .A(_2349_), .B(wData[23]), .C(wData[27]), .D(_2356_), .Y(_2680_) );
	AND2X2 AND2X2_43 ( .A(_2679_), .B(_2680_), .Y(_2681_) );
	NAND2X1 NAND2X1_407 ( .A(wData[39]), .B(_2378_), .Y(_2682_) );
	NAND2X1 NAND2X1_408 ( .A(wData[43]), .B(_2376_), .Y(_2683_) );
	NAND2X1 NAND2X1_409 ( .A(_2682_), .B(_2683_), .Y(_2684_) );
	NAND2X1 NAND2X1_410 ( .A(wData[19]), .B(_2352_), .Y(_2685_) );
	NAND2X1 NAND2X1_411 ( .A(wData[35]), .B(_2366_), .Y(_2686_) );
	NAND2X1 NAND2X1_412 ( .A(_2685_), .B(_2686_), .Y(_2687_) );
	NOR2X1 NOR2X1_230 ( .A(_2684_), .B(_2687_), .Y(_2688_) );
	NAND3X1 NAND3X1_98 ( .A(_2681_), .B(_2678_), .C(_2688_), .Y(_2689_) );
	NOR2X1 NOR2X1_231 ( .A(_2674_), .B(_2689_), .Y(_2690_) );
	AOI21X1 AOI21X1_48 ( .A(_2616_), .B(_2667_), .C(_2690_), .Y(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_3_) );
	INVX1 INVX1_250 ( .A(wSelec[55]), .Y(_2691_) );
	NOR2X1 NOR2X1_232 ( .A(wBusy_bF_buf2), .B(_2691_), .Y(_2692_) );
	INVX1 INVX1_251 ( .A(_2692_), .Y(_2693_) );
	INVX1 INVX1_252 ( .A(wSelec[65]), .Y(_2694_) );
	NAND2X1 NAND2X1_413 ( .A(wSelec[64]), .B(_2694_), .Y(_2695_) );
	INVX2 INVX2_7 ( .A(_2695_), .Y(_2696_) );
	OR2X2 OR2X2_23 ( .A(wSelec[61]), .B(wSelec[60]), .Y(_2697_) );
	INVX1 INVX1_253 ( .A(wSelec[63]), .Y(_2698_) );
	NAND2X1 NAND2X1_414 ( .A(wSelec[62]), .B(_2698_), .Y(_2699_) );
	NOR2X1 NOR2X1_233 ( .A(_2697_), .B(_2699_), .Y(_2700_) );
	AND2X2 AND2X2_44 ( .A(_2700_), .B(_2696_), .Y(_2701_) );
	AOI21X1 AOI21X1_49 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_2701_), .C(_2693_), .Y(_2702_) );
	INVX1 INVX1_254 ( .A(wSelec[61]), .Y(_2703_) );
	NAND2X1 NAND2X1_415 ( .A(wSelec[60]), .B(_2703_), .Y(_2704_) );
	OR2X2 OR2X2_24 ( .A(wSelec[62]), .B(wSelec[63]), .Y(_2705_) );
	NOR2X1 NOR2X1_234 ( .A(_2705_), .B(_2704_), .Y(_2706_) );
	NAND2X1 NAND2X1_416 ( .A(_2696_), .B(_2706_), .Y(_2707_) );
	INVX1 INVX1_255 ( .A(_2707_), .Y(_2708_) );
	INVX1 INVX1_256 ( .A(wSelec[60]), .Y(_2709_) );
	NAND2X1 NAND2X1_417 ( .A(wSelec[61]), .B(_2709_), .Y(_2710_) );
	INVX1 INVX1_257 ( .A(wSelec[62]), .Y(_2711_) );
	NAND2X1 NAND2X1_418 ( .A(wSelec[63]), .B(_2711_), .Y(_2712_) );
	NOR2X1 NOR2X1_235 ( .A(_2710_), .B(_2712_), .Y(_2713_) );
	NAND2X1 NAND2X1_419 ( .A(wSelec[64]), .B(wSelec[65]), .Y(_2714_) );
	INVX1 INVX1_258 ( .A(_2714_), .Y(_2715_) );
	NAND2X1 NAND2X1_420 ( .A(_2715_), .B(_2713_), .Y(_2716_) );
	INVX1 INVX1_259 ( .A(_2716_), .Y(_2717_) );
	AOI22X1 AOI22X1_319 ( .A(_2708_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_2717_), .Y(_2718_) );
	OR2X2 OR2X2_25 ( .A(_2704_), .B(_2705_), .Y(_2719_) );
	OR2X2 OR2X2_26 ( .A(wSelec[64]), .B(wSelec[65]), .Y(_2720_) );
	NOR2X1 NOR2X1_236 ( .A(_2720_), .B(_2719_), .Y(_2721_) );
	NOR2X1 NOR2X1_237 ( .A(_2699_), .B(_2704_), .Y(_2722_) );
	INVX1 INVX1_260 ( .A(wSelec[64]), .Y(_2723_) );
	NAND2X1 NAND2X1_421 ( .A(wSelec[65]), .B(_2723_), .Y(_2724_) );
	INVX2 INVX2_8 ( .A(_2724_), .Y(_2725_) );
	NAND2X1 NAND2X1_422 ( .A(_2725_), .B(_2722_), .Y(_2726_) );
	INVX1 INVX1_261 ( .A(_2726_), .Y(_2727_) );
	AOI22X1 AOI22X1_320 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_2721_), .C(_2727_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_2728_) );
	NAND3X1 NAND3X1_99 ( .A(_2702_), .B(_2728_), .C(_2718_), .Y(_2729_) );
	NOR2X1 NOR2X1_238 ( .A(wSelec[61]), .B(wSelec[60]), .Y(_2730_) );
	NOR2X1 NOR2X1_239 ( .A(wSelec[62]), .B(wSelec[63]), .Y(_2731_) );
	NAND2X1 NAND2X1_423 ( .A(_2730_), .B(_2731_), .Y(_2732_) );
	NOR2X1 NOR2X1_240 ( .A(_2695_), .B(_2732_), .Y(_2733_) );
	NAND2X1 NAND2X1_424 ( .A(wSelec[61]), .B(wSelec[60]), .Y(_2734_) );
	NOR3X1 NOR3X1_162 ( .A(_2705_), .B(_2734_), .C(_2695_), .Y(_2735_) );
	AOI22X1 AOI22X1_321 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_2735_), .C(_2733_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_2736_) );
	INVX1 INVX1_262 ( .A(_2720_), .Y(_2737_) );
	NOR2X1 NOR2X1_241 ( .A(_2705_), .B(_2710_), .Y(_2738_) );
	AND2X2 AND2X2_45 ( .A(_2738_), .B(_2737_), .Y(_2739_) );
	NAND2X1 NAND2X1_425 ( .A(wSelec[62]), .B(wSelec[63]), .Y(_2740_) );
	NOR3X1 NOR3X1_163 ( .A(_2714_), .B(_2734_), .C(_2740_), .Y(_2741_) );
	AOI22X1 AOI22X1_322 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_2741_), .C(_2739_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_2742_) );
	INVX1 INVX1_263 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_2743_) );
	INVX1 INVX1_264 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_2744_) );
	NOR2X1 NOR2X1_242 ( .A(_2704_), .B(_2712_), .Y(_2745_) );
	NAND2X1 NAND2X1_426 ( .A(_2715_), .B(_2745_), .Y(_2746_) );
	NOR2X1 NOR2X1_243 ( .A(_2734_), .B(_2740_), .Y(_2747_) );
	NAND2X1 NAND2X1_427 ( .A(_2747_), .B(_2725_), .Y(_2748_) );
	OAI22X1 OAI22X1_54 ( .A(_2743_), .B(_2748_), .C(_2746_), .D(_2744_), .Y(_2749_) );
	INVX1 INVX1_265 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_2750_) );
	NOR3X1 NOR3X1_164 ( .A(_2695_), .B(_2710_), .C(_2712_), .Y(_2751_) );
	NAND2X1 NAND2X1_428 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_2751_), .Y(_2752_) );
	NOR2X1 NOR2X1_244 ( .A(_2734_), .B(_2699_), .Y(_2753_) );
	NAND2X1 NAND2X1_429 ( .A(_2725_), .B(_2753_), .Y(_2754_) );
	OAI21X1 OAI21X1_70 ( .A(_2750_), .B(_2754_), .C(_2752_), .Y(_2755_) );
	NOR2X1 NOR2X1_245 ( .A(_2749_), .B(_2755_), .Y(_2756_) );
	NAND3X1 NAND3X1_100 ( .A(_2736_), .B(_2742_), .C(_2756_), .Y(_2757_) );
	INVX1 INVX1_266 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_2758_) );
	INVX1 INVX1_267 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_2759_) );
	NOR2X1 NOR2X1_246 ( .A(_2699_), .B(_2710_), .Y(_2760_) );
	NAND2X1 NAND2X1_430 ( .A(_2696_), .B(_2760_), .Y(_2761_) );
	NOR2X1 NOR2X1_247 ( .A(_2697_), .B(_2712_), .Y(_2762_) );
	NAND2X1 NAND2X1_431 ( .A(_2696_), .B(_2762_), .Y(_2763_) );
	OAI22X1 OAI22X1_55 ( .A(_2763_), .B(_2758_), .C(_2759_), .D(_2761_), .Y(_2764_) );
	INVX1 INVX1_268 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_2765_) );
	INVX1 INVX1_269 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_2766_) );
	NAND2X1 NAND2X1_432 ( .A(_2725_), .B(_2760_), .Y(_2767_) );
	NOR2X1 NOR2X1_248 ( .A(_2734_), .B(_2705_), .Y(_2768_) );
	NAND2X1 NAND2X1_433 ( .A(_2725_), .B(_2768_), .Y(_2769_) );
	OAI22X1 OAI22X1_56 ( .A(_2765_), .B(_2769_), .C(_2767_), .D(_2766_), .Y(_2770_) );
	NOR2X1 NOR2X1_249 ( .A(_2770_), .B(_2764_), .Y(_2771_) );
	NOR3X1 NOR3X1_165 ( .A(_2704_), .B(_2740_), .C(_2724_), .Y(_2772_) );
	NAND2X1 NAND2X1_434 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_2772_), .Y(_2773_) );
	NOR3X1 NOR3X1_166 ( .A(_2712_), .B(_2734_), .C(_2724_), .Y(_2774_) );
	NAND2X1 NAND2X1_435 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_2774_), .Y(_2775_) );
	NAND2X1 NAND2X1_436 ( .A(_2773_), .B(_2775_), .Y(_2776_) );
	INVX1 INVX1_270 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_2777_) );
	NAND2X1 NAND2X1_437 ( .A(_2715_), .B(_2700_), .Y(_2778_) );
	NOR3X1 NOR3X1_167 ( .A(_2710_), .B(_2712_), .C(_2724_), .Y(_2779_) );
	NAND2X1 NAND2X1_438 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_2779_), .Y(_2780_) );
	OAI21X1 OAI21X1_71 ( .A(_2777_), .B(_2778_), .C(_2780_), .Y(_2781_) );
	NOR2X1 NOR2X1_250 ( .A(_2776_), .B(_2781_), .Y(_2782_) );
	NAND2X1 NAND2X1_439 ( .A(_2771_), .B(_2782_), .Y(_2783_) );
	NOR3X1 NOR3X1_168 ( .A(_2729_), .B(_2783_), .C(_2757_), .Y(_2784_) );
	NAND2X1 NAND2X1_440 ( .A(_2696_), .B(_2753_), .Y(_2785_) );
	INVX1 INVX1_271 ( .A(_2785_), .Y(_2786_) );
	INVX1 INVX1_272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_2787_) );
	NOR3X1 NOR3X1_169 ( .A(_2697_), .B(_2720_), .C(_2699_), .Y(_2788_) );
	NAND2X1 NAND2X1_441 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_2788_), .Y(_2789_) );
	NAND2X1 NAND2X1_442 ( .A(_2737_), .B(_2760_), .Y(_2790_) );
	OAI21X1 OAI21X1_72 ( .A(_2790_), .B(_2787_), .C(_2789_), .Y(_2791_) );
	AOI21X1 AOI21X1_50 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_2786_), .C(_2791_), .Y(_2792_) );
	INVX1 INVX1_273 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_2793_) );
	INVX1 INVX1_274 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_2794_) );
	NOR2X1 NOR2X1_251 ( .A(_2740_), .B(_2697_), .Y(_2795_) );
	NAND2X1 NAND2X1_443 ( .A(_2696_), .B(_2795_), .Y(_2796_) );
	NAND2X1 NAND2X1_444 ( .A(_2737_), .B(_2722_), .Y(_2797_) );
	OAI22X1 OAI22X1_57 ( .A(_2794_), .B(_2796_), .C(_2797_), .D(_2793_), .Y(_2798_) );
	INVX1 INVX1_275 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_2799_) );
	INVX1 INVX1_276 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_2800_) );
	NAND2X1 NAND2X1_445 ( .A(_2696_), .B(_2722_), .Y(_2801_) );
	NAND2X1 NAND2X1_446 ( .A(_2737_), .B(_2768_), .Y(_2802_) );
	OAI22X1 OAI22X1_58 ( .A(_2799_), .B(_2802_), .C(_2801_), .D(_2800_), .Y(_2803_) );
	NOR2X1 NOR2X1_252 ( .A(_2798_), .B(_2803_), .Y(_2804_) );
	INVX1 INVX1_277 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_2805_) );
	NOR3X1 NOR3X1_170 ( .A(_2720_), .B(_2734_), .C(_2699_), .Y(_2806_) );
	NAND2X1 NAND2X1_447 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_2806_), .Y(_2807_) );
	OR2X2 OR2X2_27 ( .A(_2732_), .B(_2714_), .Y(_2808_) );
	OAI21X1 OAI21X1_73 ( .A(_2805_), .B(_2808_), .C(_2807_), .Y(_2809_) );
	INVX1 INVX1_278 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_2810_) );
	INVX1 INVX1_279 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_2811_) );
	NOR2X1 NOR2X1_253 ( .A(_2740_), .B(_2710_), .Y(_2812_) );
	NAND2X1 NAND2X1_448 ( .A(_2696_), .B(_2812_), .Y(_2813_) );
	NAND2X1 NAND2X1_449 ( .A(_2715_), .B(_2706_), .Y(_2814_) );
	OAI22X1 OAI22X1_59 ( .A(_2813_), .B(_2811_), .C(_2810_), .D(_2814_), .Y(_2815_) );
	NOR2X1 NOR2X1_254 ( .A(_2809_), .B(_2815_), .Y(_2816_) );
	NAND3X1 NAND3X1_101 ( .A(_2792_), .B(_2816_), .C(_2804_), .Y(_2817_) );
	NOR3X1 NOR3X1_171 ( .A(_2697_), .B(_2705_), .C(_2720_), .Y(_2818_) );
	NOR3X1 NOR3X1_172 ( .A(_2714_), .B(_2740_), .C(_2704_), .Y(_2819_) );
	AOI22X1 AOI22X1_323 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_2818_), .C(_2819_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_2820_) );
	NOR3X1 NOR3X1_173 ( .A(_2714_), .B(_2740_), .C(_2710_), .Y(_2821_) );
	NOR3X1 NOR3X1_174 ( .A(_2714_), .B(_2734_), .C(_2712_), .Y(_2822_) );
	AOI22X1 AOI22X1_324 ( .A(_2821_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_2822_), .Y(_2823_) );
	NAND2X1 NAND2X1_450 ( .A(_2820_), .B(_2823_), .Y(_2824_) );
	NOR3X1 NOR3X1_175 ( .A(_2712_), .B(_2697_), .C(_2724_), .Y(_2825_) );
	NOR3X1 NOR3X1_176 ( .A(_2704_), .B(_2712_), .C(_2724_), .Y(_2826_) );
	AOI22X1 AOI22X1_325 ( .A(_2825_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_2826_), .Y(_2827_) );
	NOR3X1 NOR3X1_177 ( .A(_2695_), .B(_2740_), .C(_2704_), .Y(_2828_) );
	NOR3X1 NOR3X1_178 ( .A(_2734_), .B(_2740_), .C(_2695_), .Y(_2829_) );
	AOI22X1 AOI22X1_326 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_2829_), .C(_2828_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_2830_) );
	NAND2X1 NAND2X1_451 ( .A(_2830_), .B(_2827_), .Y(_2831_) );
	NOR2X1 NOR2X1_255 ( .A(_2824_), .B(_2831_), .Y(_2832_) );
	NOR3X1 NOR3X1_179 ( .A(_2720_), .B(_2740_), .C(_2704_), .Y(_2833_) );
	NOR3X1 NOR3X1_180 ( .A(_2720_), .B(_2740_), .C(_2710_), .Y(_2834_) );
	AOI22X1 AOI22X1_327 ( .A(_2833_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_2834_), .Y(_2835_) );
	NOR3X1 NOR3X1_181 ( .A(_2720_), .B(_2734_), .C(_2712_), .Y(_2836_) );
	NOR3X1 NOR3X1_182 ( .A(_2695_), .B(_2705_), .C(_2710_), .Y(_2837_) );
	AOI22X1 AOI22X1_328 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_2836_), .C(_2837_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_2838_) );
	NAND2X1 NAND2X1_452 ( .A(_2835_), .B(_2838_), .Y(_2839_) );
	NOR3X1 NOR3X1_183 ( .A(_2734_), .B(_2740_), .C(_2720_), .Y(_2840_) );
	NOR3X1 NOR3X1_184 ( .A(_2710_), .B(_2705_), .C(_2724_), .Y(_2841_) );
	AOI22X1 AOI22X1_329 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_2840_), .C(_2841_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_2842_) );
	NOR3X1 NOR3X1_185 ( .A(_2697_), .B(_2705_), .C(_2724_), .Y(_2843_) );
	NOR3X1 NOR3X1_186 ( .A(_2697_), .B(_2740_), .C(_2724_), .Y(_2844_) );
	AOI22X1 AOI22X1_330 ( .A(_2843_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_2844_), .Y(_2845_) );
	NAND2X1 NAND2X1_453 ( .A(_2845_), .B(_2842_), .Y(_2846_) );
	NOR2X1 NOR2X1_256 ( .A(_2839_), .B(_2846_), .Y(_2847_) );
	NAND2X1 NAND2X1_454 ( .A(_2847_), .B(_2832_), .Y(_2848_) );
	NOR3X1 NOR3X1_187 ( .A(_2695_), .B(_2734_), .C(_2712_), .Y(_2849_) );
	NOR3X1 NOR3X1_188 ( .A(_2705_), .B(_2714_), .C(_2710_), .Y(_2850_) );
	AOI22X1 AOI22X1_331 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_2850_), .C(_2849_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_2851_) );
	NOR3X1 NOR3X1_189 ( .A(_2699_), .B(_2697_), .C(_2724_), .Y(_2852_) );
	NOR3X1 NOR3X1_190 ( .A(_2710_), .B(_2740_), .C(_2724_), .Y(_2853_) );
	AOI22X1 AOI22X1_332 ( .A(_2852_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_2853_), .Y(_2854_) );
	NAND2X1 NAND2X1_455 ( .A(_2851_), .B(_2854_), .Y(_2855_) );
	NOR3X1 NOR3X1_191 ( .A(_2695_), .B(_2704_), .C(_2712_), .Y(_2856_) );
	NAND2X1 NAND2X1_456 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_2856_), .Y(_2857_) );
	NOR3X1 NOR3X1_192 ( .A(_2714_), .B(_2734_), .C(_2699_), .Y(_2858_) );
	NAND2X1 NAND2X1_457 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_2858_), .Y(_2859_) );
	NOR3X1 NOR3X1_193 ( .A(_2697_), .B(_2740_), .C(_2720_), .Y(_2860_) );
	NOR3X1 NOR3X1_194 ( .A(_2697_), .B(_2714_), .C(_2712_), .Y(_2861_) );
	AOI22X1 AOI22X1_333 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_2860_), .C(_2861_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_2862_) );
	NAND3X1 NAND3X1_102 ( .A(_2857_), .B(_2859_), .C(_2862_), .Y(_2863_) );
	NOR2X1 NOR2X1_257 ( .A(_2863_), .B(_2855_), .Y(_2864_) );
	NOR3X1 NOR3X1_195 ( .A(_2697_), .B(_2720_), .C(_2712_), .Y(_2865_) );
	NOR3X1 NOR3X1_196 ( .A(_2699_), .B(_2714_), .C(_2704_), .Y(_2866_) );
	AOI22X1 AOI22X1_334 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_2865_), .C(_2866_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_2867_) );
	NOR3X1 NOR3X1_197 ( .A(_2699_), .B(_2714_), .C(_2710_), .Y(_2868_) );
	NAND2X1 NAND2X1_458 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_2868_), .Y(_2869_) );
	NOR3X1 NOR3X1_198 ( .A(_2704_), .B(_2705_), .C(_2724_), .Y(_2870_) );
	NAND2X1 NAND2X1_459 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_2870_), .Y(_2871_) );
	NAND3X1 NAND3X1_103 ( .A(_2869_), .B(_2871_), .C(_2867_), .Y(_2872_) );
	NOR3X1 NOR3X1_199 ( .A(_2704_), .B(_2720_), .C(_2712_), .Y(_2873_) );
	NOR3X1 NOR3X1_200 ( .A(_2714_), .B(_2740_), .C(_2697_), .Y(_2874_) );
	AOI22X1 AOI22X1_335 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_2874_), .C(_2873_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_2875_) );
	NOR3X1 NOR3X1_201 ( .A(_2710_), .B(_2720_), .C(_2712_), .Y(_2876_) );
	NOR3X1 NOR3X1_202 ( .A(_2714_), .B(_2734_), .C(_2705_), .Y(_2877_) );
	AOI22X1 AOI22X1_336 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_2877_), .C(_2876_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_2878_) );
	NAND2X1 NAND2X1_460 ( .A(_2875_), .B(_2878_), .Y(_2879_) );
	NOR2X1 NOR2X1_258 ( .A(_2879_), .B(_2872_), .Y(_2880_) );
	NAND2X1 NAND2X1_461 ( .A(_2864_), .B(_2880_), .Y(_2881_) );
	NOR3X1 NOR3X1_203 ( .A(_2848_), .B(_2817_), .C(_2881_), .Y(_2882_) );
	INVX1 INVX1_280 ( .A(wSelec[57]), .Y(_2883_) );
	NAND2X1 NAND2X1_462 ( .A(wSelec[56]), .B(_2883_), .Y(_2884_) );
	INVX1 INVX1_281 ( .A(wSelec[59]), .Y(_2885_) );
	NAND2X1 NAND2X1_463 ( .A(wSelec[58]), .B(_2885_), .Y(_2886_) );
	NOR2X1 NOR2X1_259 ( .A(_2884_), .B(_2886_), .Y(_2887_) );
	NOR2X1 NOR2X1_260 ( .A(wSelec[57]), .B(wSelec[56]), .Y(_2888_) );
	INVX1 INVX1_282 ( .A(_2888_), .Y(_2889_) );
	NOR2X1 NOR2X1_261 ( .A(_2886_), .B(_2889_), .Y(_2890_) );
	AOI22X1 AOI22X1_337 ( .A(wData[20]), .B(_2887_), .C(_2890_), .D(wData[16]), .Y(_2891_) );
	INVX1 INVX1_283 ( .A(wSelec[56]), .Y(_2892_) );
	NAND2X1 NAND2X1_464 ( .A(wSelec[57]), .B(_2892_), .Y(_2893_) );
	NOR2X1 NOR2X1_262 ( .A(_2893_), .B(_2886_), .Y(_2894_) );
	NAND2X1 NAND2X1_465 ( .A(wData[24]), .B(_2894_), .Y(_2895_) );
	INVX1 INVX1_284 ( .A(wSelec[58]), .Y(_2896_) );
	NAND2X1 NAND2X1_466 ( .A(_2896_), .B(_2885_), .Y(_2897_) );
	NOR2X1 NOR2X1_263 ( .A(_2884_), .B(_2897_), .Y(_2898_) );
	NAND2X1 NAND2X1_467 ( .A(wSelec[57]), .B(wSelec[56]), .Y(_2899_) );
	NOR2X1 NOR2X1_264 ( .A(_2899_), .B(_2886_), .Y(_2900_) );
	AOI22X1 AOI22X1_338 ( .A(_2900_), .B(wData[28]), .C(wData[4]), .D(_2898_), .Y(_2901_) );
	NAND3X1 NAND3X1_104 ( .A(_2895_), .B(_2901_), .C(_2891_), .Y(_2902_) );
	NAND2X1 NAND2X1_468 ( .A(wSelec[59]), .B(_2896_), .Y(_2903_) );
	NOR2X1 NOR2X1_265 ( .A(_2903_), .B(_2889_), .Y(_2904_) );
	NAND2X1 NAND2X1_469 ( .A(wData[32]), .B(_2904_), .Y(_2905_) );
	NAND2X1 NAND2X1_470 ( .A(wSelec[58]), .B(wSelec[59]), .Y(_2906_) );
	NOR2X1 NOR2X1_266 ( .A(_2906_), .B(_2893_), .Y(_2907_) );
	NOR2X1 NOR2X1_267 ( .A(_2906_), .B(_2884_), .Y(_2908_) );
	AOI22X1 AOI22X1_339 ( .A(_2907_), .B(wData[56]), .C(wData[52]), .D(_2908_), .Y(_2909_) );
	NOR2X1 NOR2X1_268 ( .A(_2899_), .B(_2906_), .Y(_2910_) );
	NOR2X1 NOR2X1_269 ( .A(_2899_), .B(_2903_), .Y(_2911_) );
	AOI22X1 AOI22X1_340 ( .A(wData[60]), .B(_2910_), .C(_2911_), .D(wData[44]), .Y(_2912_) );
	NAND3X1 NAND3X1_105 ( .A(_2905_), .B(_2912_), .C(_2909_), .Y(_2913_) );
	NOR2X1 NOR2X1_270 ( .A(_2893_), .B(_2903_), .Y(_2914_) );
	NAND2X1 NAND2X1_471 ( .A(wData[40]), .B(_2914_), .Y(_2915_) );
	NOR2X1 NOR2X1_271 ( .A(_2903_), .B(_2884_), .Y(_2916_) );
	NAND2X1 NAND2X1_472 ( .A(wData[36]), .B(_2916_), .Y(_2917_) );
	NOR2X1 NOR2X1_272 ( .A(_2897_), .B(_2889_), .Y(_2918_) );
	NAND2X1 NAND2X1_473 ( .A(wData[0]), .B(_2918_), .Y(_2919_) );
	NAND3X1 NAND3X1_106 ( .A(_2915_), .B(_2917_), .C(_2919_), .Y(_2920_) );
	INVX1 INVX1_285 ( .A(wData[48]), .Y(_2921_) );
	NOR2X1 NOR2X1_273 ( .A(_2896_), .B(_2885_), .Y(_2922_) );
	NAND2X1 NAND2X1_474 ( .A(_2888_), .B(_2922_), .Y(_2923_) );
	NOR2X1 NOR2X1_274 ( .A(_2893_), .B(_2897_), .Y(_2924_) );
	NOR2X1 NOR2X1_275 ( .A(_2899_), .B(_2897_), .Y(_2925_) );
	AOI22X1 AOI22X1_341 ( .A(_2924_), .B(wData[8]), .C(wData[12]), .D(_2925_), .Y(_2926_) );
	OAI21X1 OAI21X1_74 ( .A(_2921_), .B(_2923_), .C(_2926_), .Y(_2927_) );
	OR2X2 OR2X2_28 ( .A(_2927_), .B(_2920_), .Y(_2928_) );
	NOR3X1 NOR3X1_204 ( .A(_2902_), .B(_2913_), .C(_2928_), .Y(_2929_) );
	AND2X2 AND2X2_46 ( .A(_2929_), .B(_2693_), .Y(_2930_) );
	AOI21X1 AOI21X1_51 ( .A(_2784_), .B(_2882_), .C(_2930_), .Y(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_0_) );
	INVX1 INVX1_286 ( .A(_2801_), .Y(_2931_) );
	AOI21X1 AOI21X1_52 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_2931_), .C(_2693_), .Y(_2932_) );
	AOI22X1 AOI22X1_342 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_2701_), .C(_2717_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_2933_) );
	AOI22X1 AOI22X1_343 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_2721_), .C(_2727_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_2934_) );
	NAND3X1 NAND3X1_107 ( .A(_2932_), .B(_2933_), .C(_2934_), .Y(_2935_) );
	INVX1 INVX1_287 ( .A(_2761_), .Y(_2936_) );
	AOI22X1 AOI22X1_344 ( .A(_2786_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_2936_), .Y(_2937_) );
	AOI22X1 AOI22X1_345 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_2860_), .C(_2739_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_2938_) );
	INVX1 INVX1_288 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_2939_) );
	INVX1 INVX1_289 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_2940_) );
	OAI22X1 OAI22X1_60 ( .A(_2939_), .B(_2748_), .C(_2746_), .D(_2940_), .Y(_2941_) );
	INVX1 INVX1_290 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_2942_) );
	NAND2X1 NAND2X1_475 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_2849_), .Y(_2943_) );
	OAI21X1 OAI21X1_75 ( .A(_2942_), .B(_2754_), .C(_2943_), .Y(_2944_) );
	NOR2X1 NOR2X1_276 ( .A(_2941_), .B(_2944_), .Y(_2945_) );
	NAND3X1 NAND3X1_108 ( .A(_2937_), .B(_2938_), .C(_2945_), .Y(_2946_) );
	INVX1 INVX1_291 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_2947_) );
	NAND2X1 NAND2X1_476 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_2733_), .Y(_2948_) );
	OAI21X1 OAI21X1_76 ( .A(_2947_), .B(_2763_), .C(_2948_), .Y(_2949_) );
	INVX1 INVX1_292 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_2950_) );
	INVX1 INVX1_293 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_2951_) );
	OAI22X1 OAI22X1_61 ( .A(_2950_), .B(_2769_), .C(_2767_), .D(_2951_), .Y(_2952_) );
	NOR2X1 NOR2X1_277 ( .A(_2952_), .B(_2949_), .Y(_2953_) );
	AOI22X1 AOI22X1_346 ( .A(_2853_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_2826_), .Y(_2954_) );
	AND2X2 AND2X2_47 ( .A(_2700_), .B(_2715_), .Y(_2955_) );
	AOI22X1 AOI22X1_347 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_2825_), .C(_2955_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_2956_) );
	NAND3X1 NAND3X1_109 ( .A(_2954_), .B(_2956_), .C(_2953_), .Y(_2957_) );
	NOR3X1 NOR3X1_205 ( .A(_2957_), .B(_2935_), .C(_2946_), .Y(_2958_) );
	INVX1 INVX1_294 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_2959_) );
	NAND2X1 NAND2X1_477 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_2788_), .Y(_2960_) );
	OAI21X1 OAI21X1_77 ( .A(_2790_), .B(_2959_), .C(_2960_), .Y(_2961_) );
	AOI21X1 AOI21X1_53 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_2837_), .C(_2961_), .Y(_2962_) );
	INVX1 INVX1_295 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_2963_) );
	INVX1 INVX1_296 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_2964_) );
	OAI22X1 OAI22X1_62 ( .A(_2964_), .B(_2796_), .C(_2797_), .D(_2963_), .Y(_2965_) );
	INVX1 INVX1_297 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_2966_) );
	NAND2X1 NAND2X1_478 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_2806_), .Y(_2967_) );
	OAI21X1 OAI21X1_78 ( .A(_2707_), .B(_2966_), .C(_2967_), .Y(_2968_) );
	NOR2X1 NOR2X1_278 ( .A(_2968_), .B(_2965_), .Y(_2969_) );
	INVX1 INVX1_298 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_2970_) );
	INVX1 INVX1_299 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_2971_) );
	OAI22X1 OAI22X1_63 ( .A(_2802_), .B(_2971_), .C(_2808_), .D(_2970_), .Y(_2972_) );
	INVX1 INVX1_300 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_2973_) );
	NOR2X1 NOR2X1_279 ( .A(_2973_), .B(_2813_), .Y(_2974_) );
	INVX1 INVX1_301 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_2975_) );
	NOR2X1 NOR2X1_280 ( .A(_2975_), .B(_2814_), .Y(_2976_) );
	NOR3X1 NOR3X1_206 ( .A(_2974_), .B(_2972_), .C(_2976_), .Y(_2977_) );
	NAND3X1 NAND3X1_110 ( .A(_2969_), .B(_2962_), .C(_2977_), .Y(_2978_) );
	AOI22X1 AOI22X1_348 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_2818_), .C(_2819_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_2979_) );
	AOI22X1 AOI22X1_349 ( .A(_2821_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_2822_), .Y(_2980_) );
	NAND2X1 NAND2X1_479 ( .A(_2979_), .B(_2980_), .Y(_2981_) );
	AOI22X1 AOI22X1_350 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_2829_), .C(_2828_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_2982_) );
	AOI22X1 AOI22X1_351 ( .A(_2772_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_2779_), .Y(_2983_) );
	NAND2X1 NAND2X1_480 ( .A(_2982_), .B(_2983_), .Y(_2984_) );
	NOR2X1 NOR2X1_281 ( .A(_2981_), .B(_2984_), .Y(_2985_) );
	AOI22X1 AOI22X1_352 ( .A(_2833_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_2834_), .Y(_2986_) );
	AOI22X1 AOI22X1_353 ( .A(_2735_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_2836_), .Y(_2987_) );
	NAND2X1 NAND2X1_481 ( .A(_2986_), .B(_2987_), .Y(_2988_) );
	AOI22X1 AOI22X1_354 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_2840_), .C(_2841_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_2989_) );
	AOI22X1 AOI22X1_355 ( .A(_2843_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_2844_), .Y(_2990_) );
	NAND2X1 NAND2X1_482 ( .A(_2990_), .B(_2989_), .Y(_2991_) );
	NOR2X1 NOR2X1_282 ( .A(_2988_), .B(_2991_), .Y(_2992_) );
	NAND2X1 NAND2X1_483 ( .A(_2992_), .B(_2985_), .Y(_2993_) );
	AOI22X1 AOI22X1_356 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_2850_), .C(_2751_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_2994_) );
	AOI22X1 AOI22X1_357 ( .A(_2774_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_2852_), .Y(_2995_) );
	NAND2X1 NAND2X1_484 ( .A(_2994_), .B(_2995_), .Y(_2996_) );
	AOI22X1 AOI22X1_358 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_2741_), .C(_2861_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_2997_) );
	NAND2X1 NAND2X1_485 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_2856_), .Y(_2998_) );
	NAND2X1 NAND2X1_486 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_2858_), .Y(_2999_) );
	NAND3X1 NAND3X1_111 ( .A(_2998_), .B(_2999_), .C(_2997_), .Y(_3000_) );
	NOR2X1 NOR2X1_283 ( .A(_3000_), .B(_2996_), .Y(_3001_) );
	AOI22X1 AOI22X1_359 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_2865_), .C(_2866_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_3002_) );
	NAND2X1 NAND2X1_487 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_2868_), .Y(_3003_) );
	NAND2X1 NAND2X1_488 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_2870_), .Y(_3004_) );
	NAND3X1 NAND3X1_112 ( .A(_3003_), .B(_3004_), .C(_3002_), .Y(_3005_) );
	AOI22X1 AOI22X1_360 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_2874_), .C(_2873_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_3006_) );
	AOI22X1 AOI22X1_361 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_2877_), .C(_2876_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_3007_) );
	NAND2X1 NAND2X1_489 ( .A(_3006_), .B(_3007_), .Y(_3008_) );
	NOR2X1 NOR2X1_284 ( .A(_3008_), .B(_3005_), .Y(_3009_) );
	NAND2X1 NAND2X1_490 ( .A(_3001_), .B(_3009_), .Y(_3010_) );
	NOR3X1 NOR3X1_207 ( .A(_2993_), .B(_2978_), .C(_3010_), .Y(_3011_) );
	AOI21X1 AOI21X1_54 ( .A(wData[21]), .B(_2887_), .C(_2692_), .Y(_3012_) );
	AOI22X1 AOI22X1_362 ( .A(_2890_), .B(wData[17]), .C(wData[1]), .D(_2918_), .Y(_3013_) );
	AOI22X1 AOI22X1_363 ( .A(_2911_), .B(wData[45]), .C(wData[25]), .D(_2894_), .Y(_3014_) );
	NAND3X1 NAND3X1_113 ( .A(_3012_), .B(_3014_), .C(_3013_), .Y(_3015_) );
	NAND3X1 NAND3X1_114 ( .A(wData[49]), .B(_2888_), .C(_2922_), .Y(_3016_) );
	AOI22X1 AOI22X1_364 ( .A(wData[61]), .B(_2910_), .C(_2898_), .D(wData[5]), .Y(_3017_) );
	AND2X2 AND2X2_48 ( .A(_3017_), .B(_3016_), .Y(_3018_) );
	AOI22X1 AOI22X1_365 ( .A(_2907_), .B(wData[57]), .C(wData[41]), .D(_2914_), .Y(_3019_) );
	AOI22X1 AOI22X1_366 ( .A(wData[53]), .B(_2908_), .C(_2904_), .D(wData[33]), .Y(_3020_) );
	AND2X2 AND2X2_49 ( .A(_3020_), .B(_3019_), .Y(_3021_) );
	AOI22X1 AOI22X1_367 ( .A(_2924_), .B(wData[9]), .C(wData[13]), .D(_2925_), .Y(_3022_) );
	AOI22X1 AOI22X1_368 ( .A(_2900_), .B(wData[29]), .C(wData[37]), .D(_2916_), .Y(_3023_) );
	AND2X2 AND2X2_50 ( .A(_3022_), .B(_3023_), .Y(_3024_) );
	NAND3X1 NAND3X1_115 ( .A(_3018_), .B(_3024_), .C(_3021_), .Y(_3025_) );
	NOR2X1 NOR2X1_285 ( .A(_3015_), .B(_3025_), .Y(_3026_) );
	AOI21X1 AOI21X1_55 ( .A(_2958_), .B(_3011_), .C(_3026_), .Y(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_1_) );
	AOI21X1 AOI21X1_56 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_2931_), .C(_2693_), .Y(_3027_) );
	INVX1 INVX1_302 ( .A(_2790_), .Y(_3028_) );
	AOI22X1 AOI22X1_369 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_2701_), .C(_3028_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_3029_) );
	INVX1 INVX1_303 ( .A(_2802_), .Y(_3030_) );
	AOI22X1 AOI22X1_370 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_2837_), .C(_3030_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_3031_) );
	NAND3X1 NAND3X1_116 ( .A(_3031_), .B(_3027_), .C(_3029_), .Y(_3032_) );
	AOI22X1 AOI22X1_371 ( .A(_2786_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_2936_), .Y(_3033_) );
	AOI22X1 AOI22X1_372 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_2735_), .C(_2708_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_3034_) );
	INVX1 INVX1_304 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_3035_) );
	NAND2X1 NAND2X1_491 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_2825_), .Y(_3036_) );
	OAI21X1 OAI21X1_79 ( .A(_3035_), .B(_2797_), .C(_3036_), .Y(_3037_) );
	INVX1 INVX1_305 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_3038_) );
	NAND2X1 NAND2X1_492 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_2751_), .Y(_3039_) );
	OAI21X1 OAI21X1_80 ( .A(_3038_), .B(_2754_), .C(_3039_), .Y(_3040_) );
	NOR2X1 NOR2X1_286 ( .A(_3037_), .B(_3040_), .Y(_3041_) );
	NAND3X1 NAND3X1_117 ( .A(_3033_), .B(_3034_), .C(_3041_), .Y(_3042_) );
	INVX1 INVX1_306 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_3043_) );
	NAND2X1 NAND2X1_493 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_2733_), .Y(_3044_) );
	OAI21X1 OAI21X1_81 ( .A(_3043_), .B(_2763_), .C(_3044_), .Y(_3045_) );
	INVX1 INVX1_307 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_3046_) );
	INVX1 INVX1_308 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_3047_) );
	OAI22X1 OAI22X1_64 ( .A(_3046_), .B(_2769_), .C(_2767_), .D(_3047_), .Y(_3048_) );
	NOR2X1 NOR2X1_287 ( .A(_3048_), .B(_3045_), .Y(_3049_) );
	AOI22X1 AOI22X1_373 ( .A(_2853_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_2826_), .Y(_3050_) );
	AND2X2 AND2X2_51 ( .A(_2725_), .B(_2747_), .Y(_3051_) );
	AOI22X1 AOI22X1_374 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_3051_), .C(_2955_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_3052_) );
	NAND3X1 NAND3X1_118 ( .A(_3050_), .B(_3052_), .C(_3049_), .Y(_3053_) );
	NOR3X1 NOR3X1_208 ( .A(_3053_), .B(_3032_), .C(_3042_), .Y(_3054_) );
	INVX1 INVX1_309 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_3055_) );
	NOR3X1 NOR3X1_209 ( .A(_3055_), .B(_2720_), .C(_2719_), .Y(_3056_) );
	AND2X2 AND2X2_52 ( .A(_2741_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_3057_) );
	AND2X2 AND2X2_53 ( .A(_2861_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_3058_) );
	NOR3X1 NOR3X1_210 ( .A(_3058_), .B(_3057_), .C(_3056_), .Y(_3059_) );
	INVX1 INVX1_310 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_3060_) );
	INVX1 INVX1_311 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_3061_) );
	OAI22X1 OAI22X1_65 ( .A(_3061_), .B(_2796_), .C(_2746_), .D(_3060_), .Y(_3062_) );
	INVX1 INVX1_312 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_3063_) );
	INVX1 INVX1_313 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_3064_) );
	NAND2X1 NAND2X1_494 ( .A(_2737_), .B(_2738_), .Y(_3065_) );
	OAI22X1 OAI22X1_66 ( .A(_3065_), .B(_3064_), .C(_3063_), .D(_2716_), .Y(_3066_) );
	NOR2X1 NOR2X1_288 ( .A(_3062_), .B(_3066_), .Y(_3067_) );
	INVX1 INVX1_314 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_3068_) );
	NOR3X1 NOR3X1_211 ( .A(_2697_), .B(_2714_), .C(_2705_), .Y(_3069_) );
	NAND2X1 NAND2X1_495 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_3069_), .Y(_3070_) );
	OAI21X1 OAI21X1_82 ( .A(_2726_), .B(_3068_), .C(_3070_), .Y(_3071_) );
	INVX1 INVX1_315 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_3072_) );
	INVX1 INVX1_316 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_3073_) );
	OAI22X1 OAI22X1_67 ( .A(_2813_), .B(_3073_), .C(_3072_), .D(_2814_), .Y(_3074_) );
	NOR2X1 NOR2X1_289 ( .A(_3071_), .B(_3074_), .Y(_3075_) );
	NAND3X1 NAND3X1_119 ( .A(_3059_), .B(_3075_), .C(_3067_), .Y(_3076_) );
	AOI22X1 AOI22X1_375 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_2818_), .C(_2819_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_3077_) );
	AOI22X1 AOI22X1_376 ( .A(_2821_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_2822_), .Y(_3078_) );
	NAND2X1 NAND2X1_496 ( .A(_3077_), .B(_3078_), .Y(_3079_) );
	AOI22X1 AOI22X1_377 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_2829_), .C(_2828_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_3080_) );
	AOI22X1 AOI22X1_378 ( .A(_2772_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_2779_), .Y(_3081_) );
	NAND2X1 NAND2X1_497 ( .A(_3080_), .B(_3081_), .Y(_3082_) );
	NOR2X1 NOR2X1_290 ( .A(_3079_), .B(_3082_), .Y(_3083_) );
	AOI22X1 AOI22X1_379 ( .A(_2833_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_2834_), .Y(_3084_) );
	AOI22X1 AOI22X1_380 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_2860_), .C(_2836_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_3085_) );
	NAND2X1 NAND2X1_498 ( .A(_3085_), .B(_3084_), .Y(_3086_) );
	AOI22X1 AOI22X1_381 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_2840_), .C(_2841_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_3087_) );
	AOI22X1 AOI22X1_382 ( .A(_2843_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_2844_), .Y(_3088_) );
	NAND2X1 NAND2X1_499 ( .A(_3088_), .B(_3087_), .Y(_3089_) );
	NOR2X1 NOR2X1_291 ( .A(_3086_), .B(_3089_), .Y(_3090_) );
	NAND2X1 NAND2X1_500 ( .A(_3090_), .B(_3083_), .Y(_3091_) );
	AOI22X1 AOI22X1_383 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_2850_), .C(_2849_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_3092_) );
	AOI22X1 AOI22X1_384 ( .A(_2774_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_2852_), .Y(_3093_) );
	NAND2X1 NAND2X1_501 ( .A(_3092_), .B(_3093_), .Y(_3094_) );
	AOI22X1 AOI22X1_385 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_2858_), .C(_2856_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_3095_) );
	AOI22X1 AOI22X1_386 ( .A(_2788_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_2806_), .Y(_3096_) );
	NAND2X1 NAND2X1_502 ( .A(_3096_), .B(_3095_), .Y(_3097_) );
	NOR2X1 NOR2X1_292 ( .A(_3097_), .B(_3094_), .Y(_3098_) );
	AOI22X1 AOI22X1_387 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_2865_), .C(_2866_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_3099_) );
	NAND2X1 NAND2X1_503 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_2868_), .Y(_3100_) );
	NAND2X1 NAND2X1_504 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_2870_), .Y(_3101_) );
	NAND3X1 NAND3X1_120 ( .A(_3100_), .B(_3101_), .C(_3099_), .Y(_3102_) );
	AOI22X1 AOI22X1_388 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_2874_), .C(_2873_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_3103_) );
	AOI22X1 AOI22X1_389 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_2877_), .C(_2876_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_3104_) );
	NAND2X1 NAND2X1_505 ( .A(_3103_), .B(_3104_), .Y(_3105_) );
	NOR2X1 NOR2X1_293 ( .A(_3105_), .B(_3102_), .Y(_3106_) );
	NAND2X1 NAND2X1_506 ( .A(_3098_), .B(_3106_), .Y(_3107_) );
	NOR3X1 NOR3X1_212 ( .A(_3091_), .B(_3076_), .C(_3107_), .Y(_3108_) );
	AOI22X1 AOI22X1_390 ( .A(_2914_), .B(wData[42]), .C(wData[38]), .D(_2916_), .Y(_3109_) );
	AOI22X1 AOI22X1_391 ( .A(_2911_), .B(wData[46]), .C(_2918_), .D(wData[2]), .Y(_3110_) );
	NAND2X1 NAND2X1_507 ( .A(_3109_), .B(_3110_), .Y(_3111_) );
	AOI21X1 AOI21X1_57 ( .A(wData[34]), .B(_2904_), .C(_3111_), .Y(_3112_) );
	INVX1 INVX1_317 ( .A(wData[50]), .Y(_3113_) );
	AOI22X1 AOI22X1_392 ( .A(_2924_), .B(wData[10]), .C(wData[14]), .D(_2925_), .Y(_3114_) );
	OAI21X1 OAI21X1_83 ( .A(_3113_), .B(_2923_), .C(_3114_), .Y(_3115_) );
	AOI22X1 AOI22X1_393 ( .A(_2887_), .B(wData[22]), .C(wData[18]), .D(_2890_), .Y(_3116_) );
	NAND2X1 NAND2X1_508 ( .A(wData[26]), .B(_2894_), .Y(_3117_) );
	AOI22X1 AOI22X1_394 ( .A(_2900_), .B(wData[30]), .C(wData[6]), .D(_2898_), .Y(_3118_) );
	NAND3X1 NAND3X1_121 ( .A(_3117_), .B(_3118_), .C(_3116_), .Y(_3119_) );
	NOR2X1 NOR2X1_294 ( .A(_3115_), .B(_3119_), .Y(_3120_) );
	NAND2X1 NAND2X1_509 ( .A(wData[58]), .B(_2907_), .Y(_3121_) );
	NAND2X1 NAND2X1_510 ( .A(wData[54]), .B(_2908_), .Y(_3122_) );
	NAND2X1 NAND2X1_511 ( .A(_3121_), .B(_3122_), .Y(_3123_) );
	AOI21X1 AOI21X1_58 ( .A(wData[62]), .B(_2910_), .C(_3123_), .Y(_3124_) );
	NAND3X1 NAND3X1_122 ( .A(_3112_), .B(_3124_), .C(_3120_), .Y(_3125_) );
	NOR2X1 NOR2X1_295 ( .A(_2692_), .B(_3125_), .Y(_3126_) );
	AOI21X1 AOI21X1_59 ( .A(_3054_), .B(_3108_), .C(_3126_), .Y(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_2_) );
	AOI21X1 AOI21X1_60 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_2936_), .C(_2693_), .Y(_3127_) );
	AOI22X1 AOI22X1_395 ( .A(_2708_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_3028_), .Y(_3128_) );
	AOI22X1 AOI22X1_396 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_3030_), .C(_2786_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_3129_) );
	NAND3X1 NAND3X1_123 ( .A(_3129_), .B(_3127_), .C(_3128_), .Y(_3130_) );
	AOI22X1 AOI22X1_397 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_2735_), .C(_2733_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_3131_) );
	AOI22X1 AOI22X1_398 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_2806_), .C(_2931_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_3132_) );
	INVX1 INVX1_318 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_3133_) );
	INVX1 INVX1_319 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_3134_) );
	OAI22X1 OAI22X1_68 ( .A(_3133_), .B(_2748_), .C(_2797_), .D(_3134_), .Y(_3135_) );
	INVX1 INVX1_320 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_3136_) );
	NAND2X1 NAND2X1_512 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_2849_), .Y(_3137_) );
	OAI21X1 OAI21X1_84 ( .A(_3136_), .B(_2754_), .C(_3137_), .Y(_3138_) );
	NOR2X1 NOR2X1_296 ( .A(_3135_), .B(_3138_), .Y(_3139_) );
	NAND3X1 NAND3X1_124 ( .A(_3131_), .B(_3132_), .C(_3139_), .Y(_3140_) );
	AND2X2 AND2X2_54 ( .A(_2762_), .B(_2696_), .Y(_3141_) );
	AOI22X1 AOI22X1_399 ( .A(_2701_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_3141_), .Y(_3142_) );
	AND2X2 AND2X2_55 ( .A(_2760_), .B(_2725_), .Y(_3143_) );
	AND2X2 AND2X2_56 ( .A(_2768_), .B(_2725_), .Y(_3144_) );
	AOI22X1 AOI22X1_400 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_3144_), .C(_3143_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_3145_) );
	NAND2X1 NAND2X1_513 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_2853_), .Y(_3146_) );
	NAND2X1 NAND2X1_514 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_2826_), .Y(_3147_) );
	NAND2X1 NAND2X1_515 ( .A(_3146_), .B(_3147_), .Y(_3148_) );
	INVX1 INVX1_321 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_3149_) );
	NAND2X1 NAND2X1_516 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_2825_), .Y(_3150_) );
	OAI21X1 OAI21X1_85 ( .A(_3149_), .B(_2778_), .C(_3150_), .Y(_3151_) );
	NOR2X1 NOR2X1_297 ( .A(_3148_), .B(_3151_), .Y(_3152_) );
	NAND3X1 NAND3X1_125 ( .A(_3142_), .B(_3145_), .C(_3152_), .Y(_3153_) );
	NOR3X1 NOR3X1_213 ( .A(_3140_), .B(_3130_), .C(_3153_), .Y(_3154_) );
	INVX1 INVX1_322 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_3155_) );
	NAND2X1 NAND2X1_517 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_2741_), .Y(_3156_) );
	OAI21X1 OAI21X1_86 ( .A(_2746_), .B(_3155_), .C(_3156_), .Y(_3157_) );
	AOI21X1 AOI21X1_61 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_2721_), .C(_3157_), .Y(_3158_) );
	INVX1 INVX1_323 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_3159_) );
	INVX1 INVX1_324 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_3160_) );
	OAI22X1 OAI22X1_69 ( .A(_3065_), .B(_3160_), .C(_3159_), .D(_2716_), .Y(_3161_) );
	INVX1 INVX1_325 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_3162_) );
	NAND2X1 NAND2X1_518 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_2861_), .Y(_3163_) );
	OAI21X1 OAI21X1_87 ( .A(_2726_), .B(_3162_), .C(_3163_), .Y(_3164_) );
	NOR2X1 NOR2X1_298 ( .A(_3164_), .B(_3161_), .Y(_3165_) );
	INVX1 INVX1_326 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_3166_) );
	INVX1 INVX1_327 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_3167_) );
	OAI22X1 OAI22X1_70 ( .A(_2813_), .B(_3167_), .C(_3166_), .D(_2814_), .Y(_3168_) );
	INVX1 INVX1_328 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_3169_) );
	NAND2X1 NAND2X1_519 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_2860_), .Y(_3170_) );
	OAI21X1 OAI21X1_88 ( .A(_3169_), .B(_2796_), .C(_3170_), .Y(_3171_) );
	NOR2X1 NOR2X1_299 ( .A(_3171_), .B(_3168_), .Y(_3172_) );
	NAND3X1 NAND3X1_126 ( .A(_3158_), .B(_3172_), .C(_3165_), .Y(_3173_) );
	AOI22X1 AOI22X1_401 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_2818_), .C(_2819_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_3174_) );
	AOI22X1 AOI22X1_402 ( .A(_2821_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_2822_), .Y(_3175_) );
	NAND2X1 NAND2X1_520 ( .A(_3174_), .B(_3175_), .Y(_3176_) );
	AOI22X1 AOI22X1_403 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_2829_), .C(_2828_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_3177_) );
	AOI22X1 AOI22X1_404 ( .A(_2772_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_2779_), .Y(_3178_) );
	NAND2X1 NAND2X1_521 ( .A(_3177_), .B(_3178_), .Y(_3179_) );
	NOR2X1 NOR2X1_300 ( .A(_3176_), .B(_3179_), .Y(_3180_) );
	AOI22X1 AOI22X1_405 ( .A(_2833_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_2834_), .Y(_3181_) );
	AOI22X1 AOI22X1_406 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_3069_), .C(_2836_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_3182_) );
	NAND2X1 NAND2X1_522 ( .A(_3182_), .B(_3181_), .Y(_3183_) );
	AOI22X1 AOI22X1_407 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_2840_), .C(_2841_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_3184_) );
	AOI22X1 AOI22X1_408 ( .A(_2843_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_2844_), .Y(_3185_) );
	NAND2X1 NAND2X1_523 ( .A(_3185_), .B(_3184_), .Y(_3186_) );
	NOR2X1 NOR2X1_301 ( .A(_3183_), .B(_3186_), .Y(_3187_) );
	NAND2X1 NAND2X1_524 ( .A(_3187_), .B(_3180_), .Y(_3188_) );
	AOI22X1 AOI22X1_409 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_2850_), .C(_2751_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_3189_) );
	AOI22X1 AOI22X1_410 ( .A(_2774_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_2852_), .Y(_3190_) );
	NAND2X1 NAND2X1_525 ( .A(_3189_), .B(_3190_), .Y(_3191_) );
	AOI22X1 AOI22X1_411 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_2858_), .C(_2856_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_3192_) );
	AOI22X1 AOI22X1_412 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_2788_), .C(_2837_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_3193_) );
	NAND2X1 NAND2X1_526 ( .A(_3193_), .B(_3192_), .Y(_3194_) );
	NOR2X1 NOR2X1_302 ( .A(_3194_), .B(_3191_), .Y(_3195_) );
	AOI22X1 AOI22X1_413 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_2865_), .C(_2866_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_3196_) );
	NAND2X1 NAND2X1_527 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_2868_), .Y(_3197_) );
	NAND2X1 NAND2X1_528 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_2870_), .Y(_3198_) );
	NAND3X1 NAND3X1_127 ( .A(_3197_), .B(_3198_), .C(_3196_), .Y(_3199_) );
	AOI22X1 AOI22X1_414 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_2874_), .C(_2873_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_3200_) );
	AOI22X1 AOI22X1_415 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_2877_), .C(_2876_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_3201_) );
	NAND2X1 NAND2X1_529 ( .A(_3200_), .B(_3201_), .Y(_3202_) );
	NOR2X1 NOR2X1_303 ( .A(_3202_), .B(_3199_), .Y(_3203_) );
	NAND2X1 NAND2X1_530 ( .A(_3195_), .B(_3203_), .Y(_3204_) );
	NOR3X1 NOR3X1_214 ( .A(_3188_), .B(_3173_), .C(_3204_), .Y(_3205_) );
	NAND2X1 NAND2X1_531 ( .A(wData[59]), .B(_2907_), .Y(_3206_) );
	OAI21X1 OAI21X1_89 ( .A(_2691_), .B(wBusy_bF_buf1), .C(_3206_), .Y(_3207_) );
	NAND2X1 NAND2X1_532 ( .A(wData[7]), .B(_2898_), .Y(_3208_) );
	NAND2X1 NAND2X1_533 ( .A(wData[55]), .B(_2908_), .Y(_3209_) );
	AOI22X1 AOI22X1_416 ( .A(wData[63]), .B(_2910_), .C(_2900_), .D(wData[31]), .Y(_3210_) );
	NAND3X1 NAND3X1_128 ( .A(_3208_), .B(_3209_), .C(_3210_), .Y(_3211_) );
	OR2X2 OR2X2_29 ( .A(_3211_), .B(_3207_), .Y(_3212_) );
	INVX1 INVX1_329 ( .A(wData[51]), .Y(_3213_) );
	NAND2X1 NAND2X1_534 ( .A(wData[47]), .B(_2911_), .Y(_3214_) );
	OAI21X1 OAI21X1_90 ( .A(_3213_), .B(_2923_), .C(_3214_), .Y(_3215_) );
	AOI21X1 AOI21X1_62 ( .A(wData[3]), .B(_2918_), .C(_3215_), .Y(_3216_) );
	AOI22X1 AOI22X1_417 ( .A(_2924_), .B(wData[11]), .C(wData[15]), .D(_2925_), .Y(_3217_) );
	AOI22X1 AOI22X1_418 ( .A(_2887_), .B(wData[23]), .C(wData[27]), .D(_2894_), .Y(_3218_) );
	AND2X2 AND2X2_57 ( .A(_3217_), .B(_3218_), .Y(_3219_) );
	NAND2X1 NAND2X1_535 ( .A(wData[39]), .B(_2916_), .Y(_3220_) );
	NAND2X1 NAND2X1_536 ( .A(wData[43]), .B(_2914_), .Y(_3221_) );
	NAND2X1 NAND2X1_537 ( .A(_3220_), .B(_3221_), .Y(_3222_) );
	NAND2X1 NAND2X1_538 ( .A(wData[19]), .B(_2890_), .Y(_3223_) );
	NAND2X1 NAND2X1_539 ( .A(wData[35]), .B(_2904_), .Y(_3224_) );
	NAND2X1 NAND2X1_540 ( .A(_3223_), .B(_3224_), .Y(_3225_) );
	NOR2X1 NOR2X1_304 ( .A(_3222_), .B(_3225_), .Y(_3226_) );
	NAND3X1 NAND3X1_129 ( .A(_3219_), .B(_3216_), .C(_3226_), .Y(_3227_) );
	NOR2X1 NOR2X1_305 ( .A(_3212_), .B(_3227_), .Y(_3228_) );
	AOI21X1 AOI21X1_63 ( .A(_3154_), .B(_3205_), .C(_3228_), .Y(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_3_) );
	INVX1 INVX1_330 ( .A(wSelec[66]), .Y(_3229_) );
	NOR2X1 NOR2X1_306 ( .A(wBusy_bF_buf0), .B(_3229_), .Y(_3230_) );
	INVX1 INVX1_331 ( .A(_3230_), .Y(_3231_) );
	INVX1 INVX1_332 ( .A(wSelec[76]), .Y(_3232_) );
	NAND2X1 NAND2X1_541 ( .A(wSelec[75]), .B(_3232_), .Y(_3233_) );
	INVX2 INVX2_9 ( .A(_3233_), .Y(_3234_) );
	OR2X2 OR2X2_30 ( .A(wSelec[72]), .B(wSelec[71]), .Y(_3235_) );
	INVX1 INVX1_333 ( .A(wSelec[74]), .Y(_3236_) );
	NAND2X1 NAND2X1_542 ( .A(wSelec[73]), .B(_3236_), .Y(_3237_) );
	NOR2X1 NOR2X1_307 ( .A(_3235_), .B(_3237_), .Y(_3238_) );
	AND2X2 AND2X2_58 ( .A(_3238_), .B(_3234_), .Y(_3239_) );
	AOI21X1 AOI21X1_64 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_3239_), .C(_3231_), .Y(_3240_) );
	INVX1 INVX1_334 ( .A(wSelec[72]), .Y(_3241_) );
	NAND2X1 NAND2X1_543 ( .A(wSelec[71]), .B(_3241_), .Y(_3242_) );
	OR2X2 OR2X2_31 ( .A(wSelec[73]), .B(wSelec[74]), .Y(_3243_) );
	NOR2X1 NOR2X1_308 ( .A(_3243_), .B(_3242_), .Y(_3244_) );
	NAND2X1 NAND2X1_544 ( .A(_3234_), .B(_3244_), .Y(_3245_) );
	INVX1 INVX1_335 ( .A(_3245_), .Y(_3246_) );
	INVX1 INVX1_336 ( .A(wSelec[71]), .Y(_3247_) );
	NAND2X1 NAND2X1_545 ( .A(wSelec[72]), .B(_3247_), .Y(_3248_) );
	INVX1 INVX1_337 ( .A(wSelec[73]), .Y(_3249_) );
	NAND2X1 NAND2X1_546 ( .A(wSelec[74]), .B(_3249_), .Y(_3250_) );
	NOR2X1 NOR2X1_309 ( .A(_3248_), .B(_3250_), .Y(_3251_) );
	NAND2X1 NAND2X1_547 ( .A(wSelec[75]), .B(wSelec[76]), .Y(_3252_) );
	INVX1 INVX1_338 ( .A(_3252_), .Y(_3253_) );
	NAND2X1 NAND2X1_548 ( .A(_3253_), .B(_3251_), .Y(_3254_) );
	INVX1 INVX1_339 ( .A(_3254_), .Y(_3255_) );
	AOI22X1 AOI22X1_419 ( .A(_3246_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_3255_), .Y(_3256_) );
	OR2X2 OR2X2_32 ( .A(_3242_), .B(_3243_), .Y(_3257_) );
	OR2X2 OR2X2_33 ( .A(wSelec[75]), .B(wSelec[76]), .Y(_3258_) );
	NOR2X1 NOR2X1_310 ( .A(_3258_), .B(_3257_), .Y(_3259_) );
	NOR2X1 NOR2X1_311 ( .A(_3237_), .B(_3242_), .Y(_3260_) );
	INVX1 INVX1_340 ( .A(wSelec[75]), .Y(_3261_) );
	NAND2X1 NAND2X1_549 ( .A(wSelec[76]), .B(_3261_), .Y(_3262_) );
	INVX2 INVX2_10 ( .A(_3262_), .Y(_3263_) );
	NAND2X1 NAND2X1_550 ( .A(_3263_), .B(_3260_), .Y(_3264_) );
	INVX1 INVX1_341 ( .A(_3264_), .Y(_3265_) );
	AOI22X1 AOI22X1_420 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_3259_), .C(_3265_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_3266_) );
	NAND3X1 NAND3X1_130 ( .A(_3240_), .B(_3266_), .C(_3256_), .Y(_3267_) );
	NOR2X1 NOR2X1_312 ( .A(wSelec[72]), .B(wSelec[71]), .Y(_3268_) );
	NOR2X1 NOR2X1_313 ( .A(wSelec[73]), .B(wSelec[74]), .Y(_3269_) );
	NAND2X1 NAND2X1_551 ( .A(_3268_), .B(_3269_), .Y(_3270_) );
	NOR2X1 NOR2X1_314 ( .A(_3233_), .B(_3270_), .Y(_3271_) );
	NAND2X1 NAND2X1_552 ( .A(wSelec[72]), .B(wSelec[71]), .Y(_3272_) );
	NOR3X1 NOR3X1_215 ( .A(_3243_), .B(_3272_), .C(_3233_), .Y(_3273_) );
	AOI22X1 AOI22X1_421 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_3273_), .C(_3271_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_3274_) );
	INVX1 INVX1_342 ( .A(_3258_), .Y(_3275_) );
	NOR2X1 NOR2X1_315 ( .A(_3243_), .B(_3248_), .Y(_3276_) );
	AND2X2 AND2X2_59 ( .A(_3276_), .B(_3275_), .Y(_3277_) );
	NAND2X1 NAND2X1_553 ( .A(wSelec[73]), .B(wSelec[74]), .Y(_3278_) );
	NOR3X1 NOR3X1_216 ( .A(_3252_), .B(_3272_), .C(_3278_), .Y(_3279_) );
	AOI22X1 AOI22X1_422 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_3279_), .C(_3277_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_3280_) );
	INVX1 INVX1_343 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_3281_) );
	INVX1 INVX1_344 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_3282_) );
	NOR2X1 NOR2X1_316 ( .A(_3242_), .B(_3250_), .Y(_3283_) );
	NAND2X1 NAND2X1_554 ( .A(_3253_), .B(_3283_), .Y(_3284_) );
	NOR2X1 NOR2X1_317 ( .A(_3272_), .B(_3278_), .Y(_3285_) );
	NAND2X1 NAND2X1_555 ( .A(_3285_), .B(_3263_), .Y(_3286_) );
	OAI22X1 OAI22X1_71 ( .A(_3281_), .B(_3286_), .C(_3284_), .D(_3282_), .Y(_3287_) );
	INVX1 INVX1_345 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_3288_) );
	NOR3X1 NOR3X1_217 ( .A(_3233_), .B(_3248_), .C(_3250_), .Y(_3289_) );
	NAND2X1 NAND2X1_556 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_3289_), .Y(_3290_) );
	NOR2X1 NOR2X1_318 ( .A(_3272_), .B(_3237_), .Y(_3291_) );
	NAND2X1 NAND2X1_557 ( .A(_3263_), .B(_3291_), .Y(_3292_) );
	OAI21X1 OAI21X1_91 ( .A(_3288_), .B(_3292_), .C(_3290_), .Y(_3293_) );
	NOR2X1 NOR2X1_319 ( .A(_3287_), .B(_3293_), .Y(_3294_) );
	NAND3X1 NAND3X1_131 ( .A(_3274_), .B(_3280_), .C(_3294_), .Y(_3295_) );
	INVX1 INVX1_346 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_3296_) );
	INVX1 INVX1_347 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_3297_) );
	NOR2X1 NOR2X1_320 ( .A(_3237_), .B(_3248_), .Y(_3298_) );
	NAND2X1 NAND2X1_558 ( .A(_3234_), .B(_3298_), .Y(_3299_) );
	NOR2X1 NOR2X1_321 ( .A(_3235_), .B(_3250_), .Y(_3300_) );
	NAND2X1 NAND2X1_559 ( .A(_3234_), .B(_3300_), .Y(_3301_) );
	OAI22X1 OAI22X1_72 ( .A(_3301_), .B(_3296_), .C(_3297_), .D(_3299_), .Y(_3302_) );
	INVX1 INVX1_348 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_3303_) );
	INVX1 INVX1_349 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_3304_) );
	NAND2X1 NAND2X1_560 ( .A(_3263_), .B(_3298_), .Y(_3305_) );
	NOR2X1 NOR2X1_322 ( .A(_3272_), .B(_3243_), .Y(_3306_) );
	NAND2X1 NAND2X1_561 ( .A(_3263_), .B(_3306_), .Y(_3307_) );
	OAI22X1 OAI22X1_73 ( .A(_3303_), .B(_3307_), .C(_3305_), .D(_3304_), .Y(_3308_) );
	NOR2X1 NOR2X1_323 ( .A(_3308_), .B(_3302_), .Y(_3309_) );
	NOR3X1 NOR3X1_218 ( .A(_3242_), .B(_3278_), .C(_3262_), .Y(_3310_) );
	NAND2X1 NAND2X1_562 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_3310_), .Y(_3311_) );
	NOR3X1 NOR3X1_219 ( .A(_3250_), .B(_3272_), .C(_3262_), .Y(_3312_) );
	NAND2X1 NAND2X1_563 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_3312_), .Y(_3313_) );
	NAND2X1 NAND2X1_564 ( .A(_3311_), .B(_3313_), .Y(_3314_) );
	INVX1 INVX1_350 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_3315_) );
	NAND2X1 NAND2X1_565 ( .A(_3253_), .B(_3238_), .Y(_3316_) );
	NOR3X1 NOR3X1_220 ( .A(_3248_), .B(_3250_), .C(_3262_), .Y(_3317_) );
	NAND2X1 NAND2X1_566 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_3317_), .Y(_3318_) );
	OAI21X1 OAI21X1_92 ( .A(_3315_), .B(_3316_), .C(_3318_), .Y(_3319_) );
	NOR2X1 NOR2X1_324 ( .A(_3314_), .B(_3319_), .Y(_3320_) );
	NAND2X1 NAND2X1_567 ( .A(_3309_), .B(_3320_), .Y(_3321_) );
	NOR3X1 NOR3X1_221 ( .A(_3267_), .B(_3321_), .C(_3295_), .Y(_3322_) );
	NAND2X1 NAND2X1_568 ( .A(_3234_), .B(_3291_), .Y(_3323_) );
	INVX1 INVX1_351 ( .A(_3323_), .Y(_3324_) );
	INVX1 INVX1_352 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_3325_) );
	NOR3X1 NOR3X1_222 ( .A(_3235_), .B(_3258_), .C(_3237_), .Y(_3326_) );
	NAND2X1 NAND2X1_569 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_3326_), .Y(_3327_) );
	NAND2X1 NAND2X1_570 ( .A(_3275_), .B(_3298_), .Y(_3328_) );
	OAI21X1 OAI21X1_93 ( .A(_3328_), .B(_3325_), .C(_3327_), .Y(_3329_) );
	AOI21X1 AOI21X1_65 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_3324_), .C(_3329_), .Y(_3330_) );
	INVX1 INVX1_353 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_3331_) );
	INVX1 INVX1_354 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_3332_) );
	NOR2X1 NOR2X1_325 ( .A(_3278_), .B(_3235_), .Y(_3333_) );
	NAND2X1 NAND2X1_571 ( .A(_3234_), .B(_3333_), .Y(_3334_) );
	NAND2X1 NAND2X1_572 ( .A(_3275_), .B(_3260_), .Y(_3335_) );
	OAI22X1 OAI22X1_74 ( .A(_3332_), .B(_3334_), .C(_3335_), .D(_3331_), .Y(_3336_) );
	INVX1 INVX1_355 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_3337_) );
	INVX1 INVX1_356 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_3338_) );
	NAND2X1 NAND2X1_573 ( .A(_3234_), .B(_3260_), .Y(_3339_) );
	NAND2X1 NAND2X1_574 ( .A(_3275_), .B(_3306_), .Y(_3340_) );
	OAI22X1 OAI22X1_75 ( .A(_3337_), .B(_3340_), .C(_3339_), .D(_3338_), .Y(_3341_) );
	NOR2X1 NOR2X1_326 ( .A(_3336_), .B(_3341_), .Y(_3342_) );
	INVX1 INVX1_357 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_3343_) );
	NOR3X1 NOR3X1_223 ( .A(_3258_), .B(_3272_), .C(_3237_), .Y(_3344_) );
	NAND2X1 NAND2X1_575 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_3344_), .Y(_3345_) );
	OR2X2 OR2X2_34 ( .A(_3270_), .B(_3252_), .Y(_3346_) );
	OAI21X1 OAI21X1_94 ( .A(_3343_), .B(_3346_), .C(_3345_), .Y(_3347_) );
	INVX1 INVX1_358 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_3348_) );
	INVX1 INVX1_359 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_3349_) );
	NOR2X1 NOR2X1_327 ( .A(_3278_), .B(_3248_), .Y(_3350_) );
	NAND2X1 NAND2X1_576 ( .A(_3234_), .B(_3350_), .Y(_3351_) );
	NAND2X1 NAND2X1_577 ( .A(_3253_), .B(_3244_), .Y(_3352_) );
	OAI22X1 OAI22X1_76 ( .A(_3351_), .B(_3349_), .C(_3348_), .D(_3352_), .Y(_3353_) );
	NOR2X1 NOR2X1_328 ( .A(_3347_), .B(_3353_), .Y(_3354_) );
	NAND3X1 NAND3X1_132 ( .A(_3330_), .B(_3354_), .C(_3342_), .Y(_3355_) );
	NOR3X1 NOR3X1_224 ( .A(_3235_), .B(_3243_), .C(_3258_), .Y(_3356_) );
	NOR3X1 NOR3X1_225 ( .A(_3252_), .B(_3278_), .C(_3242_), .Y(_3357_) );
	AOI22X1 AOI22X1_423 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_3356_), .C(_3357_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_3358_) );
	NOR3X1 NOR3X1_226 ( .A(_3252_), .B(_3278_), .C(_3248_), .Y(_3359_) );
	NOR3X1 NOR3X1_227 ( .A(_3252_), .B(_3272_), .C(_3250_), .Y(_3360_) );
	AOI22X1 AOI22X1_424 ( .A(_3359_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_3360_), .Y(_3361_) );
	NAND2X1 NAND2X1_578 ( .A(_3358_), .B(_3361_), .Y(_3362_) );
	NOR3X1 NOR3X1_228 ( .A(_3250_), .B(_3235_), .C(_3262_), .Y(_3363_) );
	NOR3X1 NOR3X1_229 ( .A(_3242_), .B(_3250_), .C(_3262_), .Y(_3364_) );
	AOI22X1 AOI22X1_425 ( .A(_3363_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_3364_), .Y(_3365_) );
	NOR3X1 NOR3X1_230 ( .A(_3233_), .B(_3278_), .C(_3242_), .Y(_3366_) );
	NOR3X1 NOR3X1_231 ( .A(_3272_), .B(_3278_), .C(_3233_), .Y(_3367_) );
	AOI22X1 AOI22X1_426 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_3367_), .C(_3366_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_3368_) );
	NAND2X1 NAND2X1_579 ( .A(_3368_), .B(_3365_), .Y(_3369_) );
	NOR2X1 NOR2X1_329 ( .A(_3362_), .B(_3369_), .Y(_3370_) );
	NOR3X1 NOR3X1_232 ( .A(_3258_), .B(_3278_), .C(_3242_), .Y(_3371_) );
	NOR3X1 NOR3X1_233 ( .A(_3258_), .B(_3278_), .C(_3248_), .Y(_3372_) );
	AOI22X1 AOI22X1_427 ( .A(_3371_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_3372_), .Y(_3373_) );
	NOR3X1 NOR3X1_234 ( .A(_3258_), .B(_3272_), .C(_3250_), .Y(_3374_) );
	NOR3X1 NOR3X1_235 ( .A(_3233_), .B(_3243_), .C(_3248_), .Y(_3375_) );
	AOI22X1 AOI22X1_428 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_3374_), .C(_3375_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_3376_) );
	NAND2X1 NAND2X1_580 ( .A(_3373_), .B(_3376_), .Y(_3377_) );
	NOR3X1 NOR3X1_236 ( .A(_3272_), .B(_3278_), .C(_3258_), .Y(_3378_) );
	NOR3X1 NOR3X1_237 ( .A(_3248_), .B(_3243_), .C(_3262_), .Y(_3379_) );
	AOI22X1 AOI22X1_429 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_3378_), .C(_3379_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_3380_) );
	NOR3X1 NOR3X1_238 ( .A(_3235_), .B(_3243_), .C(_3262_), .Y(_3381_) );
	NOR3X1 NOR3X1_239 ( .A(_3235_), .B(_3278_), .C(_3262_), .Y(_3382_) );
	AOI22X1 AOI22X1_430 ( .A(_3381_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_3382_), .Y(_3383_) );
	NAND2X1 NAND2X1_581 ( .A(_3383_), .B(_3380_), .Y(_3384_) );
	NOR2X1 NOR2X1_330 ( .A(_3377_), .B(_3384_), .Y(_3385_) );
	NAND2X1 NAND2X1_582 ( .A(_3385_), .B(_3370_), .Y(_3386_) );
	NOR3X1 NOR3X1_240 ( .A(_3233_), .B(_3272_), .C(_3250_), .Y(_3387_) );
	NOR3X1 NOR3X1_241 ( .A(_3243_), .B(_3252_), .C(_3248_), .Y(_3388_) );
	AOI22X1 AOI22X1_431 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_3388_), .C(_3387_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_3389_) );
	NOR3X1 NOR3X1_242 ( .A(_3237_), .B(_3235_), .C(_3262_), .Y(_3390_) );
	NOR3X1 NOR3X1_243 ( .A(_3248_), .B(_3278_), .C(_3262_), .Y(_3391_) );
	AOI22X1 AOI22X1_432 ( .A(_3390_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_3391_), .Y(_3392_) );
	NAND2X1 NAND2X1_583 ( .A(_3389_), .B(_3392_), .Y(_3393_) );
	NOR3X1 NOR3X1_244 ( .A(_3233_), .B(_3242_), .C(_3250_), .Y(_3394_) );
	NAND2X1 NAND2X1_584 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_3394_), .Y(_3395_) );
	NOR3X1 NOR3X1_245 ( .A(_3252_), .B(_3272_), .C(_3237_), .Y(_3396_) );
	NAND2X1 NAND2X1_585 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_3396_), .Y(_3397_) );
	NOR3X1 NOR3X1_246 ( .A(_3235_), .B(_3278_), .C(_3258_), .Y(_3398_) );
	NOR3X1 NOR3X1_247 ( .A(_3235_), .B(_3252_), .C(_3250_), .Y(_3399_) );
	AOI22X1 AOI22X1_433 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_3398_), .C(_3399_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_3400_) );
	NAND3X1 NAND3X1_133 ( .A(_3395_), .B(_3397_), .C(_3400_), .Y(_3401_) );
	NOR2X1 NOR2X1_331 ( .A(_3401_), .B(_3393_), .Y(_3402_) );
	NOR3X1 NOR3X1_248 ( .A(_3235_), .B(_3258_), .C(_3250_), .Y(_3403_) );
	NOR3X1 NOR3X1_249 ( .A(_3237_), .B(_3252_), .C(_3242_), .Y(_3404_) );
	AOI22X1 AOI22X1_434 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_3403_), .C(_3404_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_3405_) );
	NOR3X1 NOR3X1_250 ( .A(_3237_), .B(_3252_), .C(_3248_), .Y(_3406_) );
	NAND2X1 NAND2X1_586 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_3406_), .Y(_3407_) );
	NOR3X1 NOR3X1_251 ( .A(_3242_), .B(_3243_), .C(_3262_), .Y(_3408_) );
	NAND2X1 NAND2X1_587 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_3408_), .Y(_3409_) );
	NAND3X1 NAND3X1_134 ( .A(_3407_), .B(_3409_), .C(_3405_), .Y(_3410_) );
	NOR3X1 NOR3X1_252 ( .A(_3242_), .B(_3258_), .C(_3250_), .Y(_3411_) );
	NOR3X1 NOR3X1_253 ( .A(_3252_), .B(_3278_), .C(_3235_), .Y(_3412_) );
	AOI22X1 AOI22X1_435 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_3412_), .C(_3411_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_3413_) );
	NOR3X1 NOR3X1_254 ( .A(_3248_), .B(_3258_), .C(_3250_), .Y(_3414_) );
	NOR3X1 NOR3X1_255 ( .A(_3252_), .B(_3272_), .C(_3243_), .Y(_3415_) );
	AOI22X1 AOI22X1_436 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_3415_), .C(_3414_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_3416_) );
	NAND2X1 NAND2X1_588 ( .A(_3413_), .B(_3416_), .Y(_3417_) );
	NOR2X1 NOR2X1_332 ( .A(_3417_), .B(_3410_), .Y(_3418_) );
	NAND2X1 NAND2X1_589 ( .A(_3402_), .B(_3418_), .Y(_3419_) );
	NOR3X1 NOR3X1_256 ( .A(_3386_), .B(_3355_), .C(_3419_), .Y(_3420_) );
	INVX1 INVX1_360 ( .A(wSelec[68]), .Y(_3421_) );
	NAND2X1 NAND2X1_590 ( .A(wSelec[67]), .B(_3421_), .Y(_3422_) );
	INVX1 INVX1_361 ( .A(wSelec[70]), .Y(_3423_) );
	NAND2X1 NAND2X1_591 ( .A(wSelec[69]), .B(_3423_), .Y(_3424_) );
	NOR2X1 NOR2X1_333 ( .A(_3422_), .B(_3424_), .Y(_3425_) );
	NOR2X1 NOR2X1_334 ( .A(wSelec[68]), .B(wSelec[67]), .Y(_3426_) );
	INVX1 INVX1_362 ( .A(_3426_), .Y(_3427_) );
	NOR2X1 NOR2X1_335 ( .A(_3424_), .B(_3427_), .Y(_3428_) );
	AOI22X1 AOI22X1_437 ( .A(wData[20]), .B(_3425_), .C(_3428_), .D(wData[16]), .Y(_3429_) );
	INVX1 INVX1_363 ( .A(wSelec[67]), .Y(_3430_) );
	NAND2X1 NAND2X1_592 ( .A(wSelec[68]), .B(_3430_), .Y(_3431_) );
	NOR2X1 NOR2X1_336 ( .A(_3431_), .B(_3424_), .Y(_3432_) );
	NAND2X1 NAND2X1_593 ( .A(wData[24]), .B(_3432_), .Y(_3433_) );
	INVX1 INVX1_364 ( .A(wSelec[69]), .Y(_3434_) );
	NAND2X1 NAND2X1_594 ( .A(_3434_), .B(_3423_), .Y(_3435_) );
	NOR2X1 NOR2X1_337 ( .A(_3422_), .B(_3435_), .Y(_3436_) );
	NAND2X1 NAND2X1_595 ( .A(wSelec[68]), .B(wSelec[67]), .Y(_3437_) );
	NOR2X1 NOR2X1_338 ( .A(_3437_), .B(_3424_), .Y(_3438_) );
	AOI22X1 AOI22X1_438 ( .A(_3438_), .B(wData[28]), .C(wData[4]), .D(_3436_), .Y(_3439_) );
	NAND3X1 NAND3X1_135 ( .A(_3433_), .B(_3439_), .C(_3429_), .Y(_3440_) );
	NAND2X1 NAND2X1_596 ( .A(wSelec[70]), .B(_3434_), .Y(_3441_) );
	NOR2X1 NOR2X1_339 ( .A(_3441_), .B(_3427_), .Y(_3442_) );
	NAND2X1 NAND2X1_597 ( .A(wData[32]), .B(_3442_), .Y(_3443_) );
	NAND2X1 NAND2X1_598 ( .A(wSelec[69]), .B(wSelec[70]), .Y(_3444_) );
	NOR2X1 NOR2X1_340 ( .A(_3444_), .B(_3431_), .Y(_3445_) );
	NOR2X1 NOR2X1_341 ( .A(_3444_), .B(_3422_), .Y(_3446_) );
	AOI22X1 AOI22X1_439 ( .A(_3445_), .B(wData[56]), .C(wData[52]), .D(_3446_), .Y(_3447_) );
	NOR2X1 NOR2X1_342 ( .A(_3437_), .B(_3444_), .Y(_3448_) );
	NOR2X1 NOR2X1_343 ( .A(_3437_), .B(_3441_), .Y(_3449_) );
	AOI22X1 AOI22X1_440 ( .A(wData[60]), .B(_3448_), .C(_3449_), .D(wData[44]), .Y(_3450_) );
	NAND3X1 NAND3X1_136 ( .A(_3443_), .B(_3450_), .C(_3447_), .Y(_3451_) );
	NOR2X1 NOR2X1_344 ( .A(_3431_), .B(_3441_), .Y(_3452_) );
	NAND2X1 NAND2X1_599 ( .A(wData[40]), .B(_3452_), .Y(_3453_) );
	NOR2X1 NOR2X1_345 ( .A(_3441_), .B(_3422_), .Y(_3454_) );
	NAND2X1 NAND2X1_600 ( .A(wData[36]), .B(_3454_), .Y(_3455_) );
	NOR2X1 NOR2X1_346 ( .A(_3435_), .B(_3427_), .Y(_3456_) );
	NAND2X1 NAND2X1_601 ( .A(wData[0]), .B(_3456_), .Y(_3457_) );
	NAND3X1 NAND3X1_137 ( .A(_3453_), .B(_3455_), .C(_3457_), .Y(_3458_) );
	INVX1 INVX1_365 ( .A(wData[48]), .Y(_3459_) );
	NOR2X1 NOR2X1_347 ( .A(_3434_), .B(_3423_), .Y(_3460_) );
	NAND2X1 NAND2X1_602 ( .A(_3426_), .B(_3460_), .Y(_3461_) );
	NOR2X1 NOR2X1_348 ( .A(_3431_), .B(_3435_), .Y(_3462_) );
	NOR2X1 NOR2X1_349 ( .A(_3437_), .B(_3435_), .Y(_3463_) );
	AOI22X1 AOI22X1_441 ( .A(_3462_), .B(wData[8]), .C(wData[12]), .D(_3463_), .Y(_3464_) );
	OAI21X1 OAI21X1_95 ( .A(_3459_), .B(_3461_), .C(_3464_), .Y(_3465_) );
	OR2X2 OR2X2_35 ( .A(_3465_), .B(_3458_), .Y(_3466_) );
	NOR3X1 NOR3X1_257 ( .A(_3440_), .B(_3451_), .C(_3466_), .Y(_3467_) );
	AND2X2 AND2X2_60 ( .A(_3467_), .B(_3231_), .Y(_3468_) );
	AOI21X1 AOI21X1_66 ( .A(_3322_), .B(_3420_), .C(_3468_), .Y(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_0_) );
	INVX1 INVX1_366 ( .A(_3339_), .Y(_3469_) );
	AOI21X1 AOI21X1_67 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_3469_), .C(_3231_), .Y(_3470_) );
	AOI22X1 AOI22X1_442 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_3239_), .C(_3255_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_3471_) );
	AOI22X1 AOI22X1_443 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_3259_), .C(_3265_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_3472_) );
	NAND3X1 NAND3X1_138 ( .A(_3470_), .B(_3471_), .C(_3472_), .Y(_3473_) );
	INVX1 INVX1_367 ( .A(_3299_), .Y(_3474_) );
	AOI22X1 AOI22X1_444 ( .A(_3324_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_3474_), .Y(_3475_) );
	AOI22X1 AOI22X1_445 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_3398_), .C(_3277_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_3476_) );
	INVX1 INVX1_368 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_3477_) );
	INVX1 INVX1_369 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_3478_) );
	OAI22X1 OAI22X1_77 ( .A(_3477_), .B(_3286_), .C(_3284_), .D(_3478_), .Y(_3479_) );
	INVX1 INVX1_370 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_3480_) );
	NAND2X1 NAND2X1_603 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_3387_), .Y(_3481_) );
	OAI21X1 OAI21X1_96 ( .A(_3480_), .B(_3292_), .C(_3481_), .Y(_3482_) );
	NOR2X1 NOR2X1_350 ( .A(_3479_), .B(_3482_), .Y(_3483_) );
	NAND3X1 NAND3X1_139 ( .A(_3475_), .B(_3476_), .C(_3483_), .Y(_3484_) );
	INVX1 INVX1_371 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_3485_) );
	NAND2X1 NAND2X1_604 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_3271_), .Y(_3486_) );
	OAI21X1 OAI21X1_97 ( .A(_3485_), .B(_3301_), .C(_3486_), .Y(_3487_) );
	INVX1 INVX1_372 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_3488_) );
	INVX1 INVX1_373 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_3489_) );
	OAI22X1 OAI22X1_78 ( .A(_3488_), .B(_3307_), .C(_3305_), .D(_3489_), .Y(_3490_) );
	NOR2X1 NOR2X1_351 ( .A(_3490_), .B(_3487_), .Y(_3491_) );
	AOI22X1 AOI22X1_446 ( .A(_3391_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_3364_), .Y(_3492_) );
	AND2X2 AND2X2_61 ( .A(_3238_), .B(_3253_), .Y(_3493_) );
	AOI22X1 AOI22X1_447 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_3363_), .C(_3493_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_3494_) );
	NAND3X1 NAND3X1_140 ( .A(_3492_), .B(_3494_), .C(_3491_), .Y(_3495_) );
	NOR3X1 NOR3X1_258 ( .A(_3495_), .B(_3473_), .C(_3484_), .Y(_3496_) );
	INVX1 INVX1_374 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_3497_) );
	NAND2X1 NAND2X1_605 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_3326_), .Y(_3498_) );
	OAI21X1 OAI21X1_98 ( .A(_3328_), .B(_3497_), .C(_3498_), .Y(_3499_) );
	AOI21X1 AOI21X1_68 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_3375_), .C(_3499_), .Y(_3500_) );
	INVX1 INVX1_375 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_3501_) );
	INVX1 INVX1_376 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_3502_) );
	OAI22X1 OAI22X1_79 ( .A(_3502_), .B(_3334_), .C(_3335_), .D(_3501_), .Y(_3503_) );
	INVX1 INVX1_377 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_3504_) );
	NAND2X1 NAND2X1_606 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_3344_), .Y(_3505_) );
	OAI21X1 OAI21X1_99 ( .A(_3245_), .B(_3504_), .C(_3505_), .Y(_3506_) );
	NOR2X1 NOR2X1_352 ( .A(_3506_), .B(_3503_), .Y(_3507_) );
	INVX1 INVX1_378 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_3508_) );
	INVX1 INVX1_379 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_3509_) );
	OAI22X1 OAI22X1_80 ( .A(_3340_), .B(_3509_), .C(_3346_), .D(_3508_), .Y(_3510_) );
	INVX1 INVX1_380 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_3511_) );
	NOR2X1 NOR2X1_353 ( .A(_3511_), .B(_3351_), .Y(_3512_) );
	INVX1 INVX1_381 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_3513_) );
	NOR2X1 NOR2X1_354 ( .A(_3513_), .B(_3352_), .Y(_3514_) );
	NOR3X1 NOR3X1_259 ( .A(_3512_), .B(_3510_), .C(_3514_), .Y(_3515_) );
	NAND3X1 NAND3X1_141 ( .A(_3507_), .B(_3500_), .C(_3515_), .Y(_3516_) );
	AOI22X1 AOI22X1_448 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_3356_), .C(_3357_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_3517_) );
	AOI22X1 AOI22X1_449 ( .A(_3359_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_3360_), .Y(_3518_) );
	NAND2X1 NAND2X1_607 ( .A(_3517_), .B(_3518_), .Y(_3519_) );
	AOI22X1 AOI22X1_450 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_3367_), .C(_3366_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_3520_) );
	AOI22X1 AOI22X1_451 ( .A(_3310_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_3317_), .Y(_3521_) );
	NAND2X1 NAND2X1_608 ( .A(_3520_), .B(_3521_), .Y(_3522_) );
	NOR2X1 NOR2X1_355 ( .A(_3519_), .B(_3522_), .Y(_3523_) );
	AOI22X1 AOI22X1_452 ( .A(_3371_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_3372_), .Y(_3524_) );
	AOI22X1 AOI22X1_453 ( .A(_3273_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_3374_), .Y(_3525_) );
	NAND2X1 NAND2X1_609 ( .A(_3524_), .B(_3525_), .Y(_3526_) );
	AOI22X1 AOI22X1_454 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_3378_), .C(_3379_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_3527_) );
	AOI22X1 AOI22X1_455 ( .A(_3381_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_3382_), .Y(_3528_) );
	NAND2X1 NAND2X1_610 ( .A(_3528_), .B(_3527_), .Y(_3529_) );
	NOR2X1 NOR2X1_356 ( .A(_3526_), .B(_3529_), .Y(_3530_) );
	NAND2X1 NAND2X1_611 ( .A(_3530_), .B(_3523_), .Y(_3531_) );
	AOI22X1 AOI22X1_456 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_3388_), .C(_3289_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_3532_) );
	AOI22X1 AOI22X1_457 ( .A(_3312_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_3390_), .Y(_3533_) );
	NAND2X1 NAND2X1_612 ( .A(_3532_), .B(_3533_), .Y(_3534_) );
	AOI22X1 AOI22X1_458 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_3279_), .C(_3399_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_3535_) );
	NAND2X1 NAND2X1_613 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_3394_), .Y(_3536_) );
	NAND2X1 NAND2X1_614 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_3396_), .Y(_3537_) );
	NAND3X1 NAND3X1_142 ( .A(_3536_), .B(_3537_), .C(_3535_), .Y(_3538_) );
	NOR2X1 NOR2X1_357 ( .A(_3538_), .B(_3534_), .Y(_3539_) );
	AOI22X1 AOI22X1_459 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_3403_), .C(_3404_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_3540_) );
	NAND2X1 NAND2X1_615 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_3406_), .Y(_3541_) );
	NAND2X1 NAND2X1_616 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_3408_), .Y(_3542_) );
	NAND3X1 NAND3X1_143 ( .A(_3541_), .B(_3542_), .C(_3540_), .Y(_3543_) );
	AOI22X1 AOI22X1_460 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_3412_), .C(_3411_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_3544_) );
	AOI22X1 AOI22X1_461 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_3415_), .C(_3414_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_3545_) );
	NAND2X1 NAND2X1_617 ( .A(_3544_), .B(_3545_), .Y(_3546_) );
	NOR2X1 NOR2X1_358 ( .A(_3546_), .B(_3543_), .Y(_3547_) );
	NAND2X1 NAND2X1_618 ( .A(_3539_), .B(_3547_), .Y(_3548_) );
	NOR3X1 NOR3X1_260 ( .A(_3531_), .B(_3516_), .C(_3548_), .Y(_3549_) );
	AOI21X1 AOI21X1_69 ( .A(wData[21]), .B(_3425_), .C(_3230_), .Y(_3550_) );
	AOI22X1 AOI22X1_462 ( .A(_3428_), .B(wData[17]), .C(wData[1]), .D(_3456_), .Y(_3551_) );
	AOI22X1 AOI22X1_463 ( .A(_3449_), .B(wData[45]), .C(wData[25]), .D(_3432_), .Y(_3552_) );
	NAND3X1 NAND3X1_144 ( .A(_3550_), .B(_3552_), .C(_3551_), .Y(_3553_) );
	NAND3X1 NAND3X1_145 ( .A(wData[49]), .B(_3426_), .C(_3460_), .Y(_3554_) );
	AOI22X1 AOI22X1_464 ( .A(wData[61]), .B(_3448_), .C(_3436_), .D(wData[5]), .Y(_3555_) );
	AND2X2 AND2X2_62 ( .A(_3555_), .B(_3554_), .Y(_3556_) );
	AOI22X1 AOI22X1_465 ( .A(_3445_), .B(wData[57]), .C(wData[41]), .D(_3452_), .Y(_3557_) );
	AOI22X1 AOI22X1_466 ( .A(wData[53]), .B(_3446_), .C(_3442_), .D(wData[33]), .Y(_3558_) );
	AND2X2 AND2X2_63 ( .A(_3558_), .B(_3557_), .Y(_3559_) );
	AOI22X1 AOI22X1_467 ( .A(_3462_), .B(wData[9]), .C(wData[13]), .D(_3463_), .Y(_3560_) );
	AOI22X1 AOI22X1_468 ( .A(_3438_), .B(wData[29]), .C(wData[37]), .D(_3454_), .Y(_3561_) );
	AND2X2 AND2X2_64 ( .A(_3560_), .B(_3561_), .Y(_3562_) );
	NAND3X1 NAND3X1_146 ( .A(_3556_), .B(_3562_), .C(_3559_), .Y(_3563_) );
	NOR2X1 NOR2X1_359 ( .A(_3553_), .B(_3563_), .Y(_3564_) );
	AOI21X1 AOI21X1_70 ( .A(_3496_), .B(_3549_), .C(_3564_), .Y(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_1_) );
	AOI21X1 AOI21X1_71 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_3469_), .C(_3231_), .Y(_3565_) );
	INVX1 INVX1_382 ( .A(_3328_), .Y(_3566_) );
	AOI22X1 AOI22X1_469 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_3239_), .C(_3566_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_3567_) );
	INVX1 INVX1_383 ( .A(_3340_), .Y(_3568_) );
	AOI22X1 AOI22X1_470 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_3375_), .C(_3568_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_3569_) );
	NAND3X1 NAND3X1_147 ( .A(_3569_), .B(_3565_), .C(_3567_), .Y(_3570_) );
	AOI22X1 AOI22X1_471 ( .A(_3324_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_3474_), .Y(_3571_) );
	AOI22X1 AOI22X1_472 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_3273_), .C(_3246_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_3572_) );
	INVX1 INVX1_384 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_3573_) );
	NAND2X1 NAND2X1_619 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_3363_), .Y(_3574_) );
	OAI21X1 OAI21X1_100 ( .A(_3573_), .B(_3335_), .C(_3574_), .Y(_3575_) );
	INVX1 INVX1_385 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_3576_) );
	NAND2X1 NAND2X1_620 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_3289_), .Y(_3577_) );
	OAI21X1 OAI21X1_101 ( .A(_3576_), .B(_3292_), .C(_3577_), .Y(_3578_) );
	NOR2X1 NOR2X1_360 ( .A(_3575_), .B(_3578_), .Y(_3579_) );
	NAND3X1 NAND3X1_148 ( .A(_3571_), .B(_3572_), .C(_3579_), .Y(_3580_) );
	INVX1 INVX1_386 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_3581_) );
	NAND2X1 NAND2X1_621 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_3271_), .Y(_3582_) );
	OAI21X1 OAI21X1_102 ( .A(_3581_), .B(_3301_), .C(_3582_), .Y(_3583_) );
	INVX1 INVX1_387 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_3584_) );
	INVX1 INVX1_388 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_3585_) );
	OAI22X1 OAI22X1_81 ( .A(_3584_), .B(_3307_), .C(_3305_), .D(_3585_), .Y(_3586_) );
	NOR2X1 NOR2X1_361 ( .A(_3586_), .B(_3583_), .Y(_3587_) );
	AOI22X1 AOI22X1_473 ( .A(_3391_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_3364_), .Y(_3588_) );
	AND2X2 AND2X2_65 ( .A(_3263_), .B(_3285_), .Y(_3589_) );
	AOI22X1 AOI22X1_474 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_3589_), .C(_3493_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_3590_) );
	NAND3X1 NAND3X1_149 ( .A(_3588_), .B(_3590_), .C(_3587_), .Y(_3591_) );
	NOR3X1 NOR3X1_261 ( .A(_3591_), .B(_3570_), .C(_3580_), .Y(_3592_) );
	INVX1 INVX1_389 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_3593_) );
	NOR3X1 NOR3X1_262 ( .A(_3593_), .B(_3258_), .C(_3257_), .Y(_3594_) );
	AND2X2 AND2X2_66 ( .A(_3279_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_3595_) );
	AND2X2 AND2X2_67 ( .A(_3399_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_3596_) );
	NOR3X1 NOR3X1_263 ( .A(_3596_), .B(_3595_), .C(_3594_), .Y(_3597_) );
	INVX1 INVX1_390 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_3598_) );
	INVX1 INVX1_391 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_3599_) );
	OAI22X1 OAI22X1_82 ( .A(_3599_), .B(_3334_), .C(_3284_), .D(_3598_), .Y(_3600_) );
	INVX1 INVX1_392 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_3601_) );
	INVX1 INVX1_393 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_3602_) );
	NAND2X1 NAND2X1_622 ( .A(_3275_), .B(_3276_), .Y(_3603_) );
	OAI22X1 OAI22X1_83 ( .A(_3603_), .B(_3602_), .C(_3601_), .D(_3254_), .Y(_3604_) );
	NOR2X1 NOR2X1_362 ( .A(_3600_), .B(_3604_), .Y(_3605_) );
	INVX1 INVX1_394 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_3606_) );
	NOR3X1 NOR3X1_264 ( .A(_3235_), .B(_3252_), .C(_3243_), .Y(_3607_) );
	NAND2X1 NAND2X1_623 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_3607_), .Y(_3608_) );
	OAI21X1 OAI21X1_103 ( .A(_3264_), .B(_3606_), .C(_3608_), .Y(_3609_) );
	INVX1 INVX1_395 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_3610_) );
	INVX1 INVX1_396 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_3611_) );
	OAI22X1 OAI22X1_84 ( .A(_3351_), .B(_3611_), .C(_3610_), .D(_3352_), .Y(_3612_) );
	NOR2X1 NOR2X1_363 ( .A(_3609_), .B(_3612_), .Y(_3613_) );
	NAND3X1 NAND3X1_150 ( .A(_3597_), .B(_3613_), .C(_3605_), .Y(_3614_) );
	AOI22X1 AOI22X1_475 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_3356_), .C(_3357_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_3615_) );
	AOI22X1 AOI22X1_476 ( .A(_3359_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_3360_), .Y(_3616_) );
	NAND2X1 NAND2X1_624 ( .A(_3615_), .B(_3616_), .Y(_3617_) );
	AOI22X1 AOI22X1_477 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_3367_), .C(_3366_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_3618_) );
	AOI22X1 AOI22X1_478 ( .A(_3310_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_3317_), .Y(_3619_) );
	NAND2X1 NAND2X1_625 ( .A(_3618_), .B(_3619_), .Y(_3620_) );
	NOR2X1 NOR2X1_364 ( .A(_3617_), .B(_3620_), .Y(_3621_) );
	AOI22X1 AOI22X1_479 ( .A(_3371_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_3372_), .Y(_3622_) );
	AOI22X1 AOI22X1_480 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_3398_), .C(_3374_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_3623_) );
	NAND2X1 NAND2X1_626 ( .A(_3623_), .B(_3622_), .Y(_3624_) );
	AOI22X1 AOI22X1_481 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_3378_), .C(_3379_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_3625_) );
	AOI22X1 AOI22X1_482 ( .A(_3381_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_3382_), .Y(_3626_) );
	NAND2X1 NAND2X1_627 ( .A(_3626_), .B(_3625_), .Y(_3627_) );
	NOR2X1 NOR2X1_365 ( .A(_3624_), .B(_3627_), .Y(_3628_) );
	NAND2X1 NAND2X1_628 ( .A(_3628_), .B(_3621_), .Y(_3629_) );
	AOI22X1 AOI22X1_483 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_3388_), .C(_3387_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_3630_) );
	AOI22X1 AOI22X1_484 ( .A(_3312_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_3390_), .Y(_3631_) );
	NAND2X1 NAND2X1_629 ( .A(_3630_), .B(_3631_), .Y(_3632_) );
	AOI22X1 AOI22X1_485 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_3396_), .C(_3394_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_3633_) );
	AOI22X1 AOI22X1_486 ( .A(_3326_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_3344_), .Y(_3634_) );
	NAND2X1 NAND2X1_630 ( .A(_3634_), .B(_3633_), .Y(_3635_) );
	NOR2X1 NOR2X1_366 ( .A(_3635_), .B(_3632_), .Y(_3636_) );
	AOI22X1 AOI22X1_487 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_3403_), .C(_3404_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_3637_) );
	NAND2X1 NAND2X1_631 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_3406_), .Y(_3638_) );
	NAND2X1 NAND2X1_632 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_3408_), .Y(_3639_) );
	NAND3X1 NAND3X1_151 ( .A(_3638_), .B(_3639_), .C(_3637_), .Y(_3640_) );
	AOI22X1 AOI22X1_488 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_3412_), .C(_3411_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_3641_) );
	AOI22X1 AOI22X1_489 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_3415_), .C(_3414_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_3642_) );
	NAND2X1 NAND2X1_633 ( .A(_3641_), .B(_3642_), .Y(_3643_) );
	NOR2X1 NOR2X1_367 ( .A(_3643_), .B(_3640_), .Y(_3644_) );
	NAND2X1 NAND2X1_634 ( .A(_3636_), .B(_3644_), .Y(_3645_) );
	NOR3X1 NOR3X1_265 ( .A(_3629_), .B(_3614_), .C(_3645_), .Y(_3646_) );
	AOI22X1 AOI22X1_490 ( .A(_3452_), .B(wData[42]), .C(wData[38]), .D(_3454_), .Y(_3647_) );
	AOI22X1 AOI22X1_491 ( .A(_3449_), .B(wData[46]), .C(_3456_), .D(wData[2]), .Y(_3648_) );
	NAND2X1 NAND2X1_635 ( .A(_3647_), .B(_3648_), .Y(_3649_) );
	AOI21X1 AOI21X1_72 ( .A(wData[34]), .B(_3442_), .C(_3649_), .Y(_3650_) );
	INVX1 INVX1_397 ( .A(wData[50]), .Y(_3651_) );
	AOI22X1 AOI22X1_492 ( .A(_3462_), .B(wData[10]), .C(wData[14]), .D(_3463_), .Y(_3652_) );
	OAI21X1 OAI21X1_104 ( .A(_3651_), .B(_3461_), .C(_3652_), .Y(_3653_) );
	AOI22X1 AOI22X1_493 ( .A(_3425_), .B(wData[22]), .C(wData[18]), .D(_3428_), .Y(_3654_) );
	NAND2X1 NAND2X1_636 ( .A(wData[26]), .B(_3432_), .Y(_3655_) );
	AOI22X1 AOI22X1_494 ( .A(_3438_), .B(wData[30]), .C(wData[6]), .D(_3436_), .Y(_3656_) );
	NAND3X1 NAND3X1_152 ( .A(_3655_), .B(_3656_), .C(_3654_), .Y(_3657_) );
	NOR2X1 NOR2X1_368 ( .A(_3653_), .B(_3657_), .Y(_3658_) );
	NAND2X1 NAND2X1_637 ( .A(wData[58]), .B(_3445_), .Y(_3659_) );
	NAND2X1 NAND2X1_638 ( .A(wData[54]), .B(_3446_), .Y(_3660_) );
	NAND2X1 NAND2X1_639 ( .A(_3659_), .B(_3660_), .Y(_3661_) );
	AOI21X1 AOI21X1_73 ( .A(wData[62]), .B(_3448_), .C(_3661_), .Y(_3662_) );
	NAND3X1 NAND3X1_153 ( .A(_3650_), .B(_3662_), .C(_3658_), .Y(_3663_) );
	NOR2X1 NOR2X1_369 ( .A(_3230_), .B(_3663_), .Y(_3664_) );
	AOI21X1 AOI21X1_74 ( .A(_3592_), .B(_3646_), .C(_3664_), .Y(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_2_) );
	AOI21X1 AOI21X1_75 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_3474_), .C(_3231_), .Y(_3665_) );
	AOI22X1 AOI22X1_495 ( .A(_3246_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_3566_), .Y(_3666_) );
	AOI22X1 AOI22X1_496 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_3568_), .C(_3324_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_3667_) );
	NAND3X1 NAND3X1_154 ( .A(_3667_), .B(_3665_), .C(_3666_), .Y(_3668_) );
	AOI22X1 AOI22X1_497 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_3273_), .C(_3271_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_3669_) );
	AOI22X1 AOI22X1_498 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_3344_), .C(_3469_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_3670_) );
	INVX1 INVX1_398 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_3671_) );
	INVX1 INVX1_399 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_3672_) );
	OAI22X1 OAI22X1_85 ( .A(_3671_), .B(_3286_), .C(_3335_), .D(_3672_), .Y(_3673_) );
	INVX1 INVX1_400 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_3674_) );
	NAND2X1 NAND2X1_640 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_3387_), .Y(_3675_) );
	OAI21X1 OAI21X1_105 ( .A(_3674_), .B(_3292_), .C(_3675_), .Y(_3676_) );
	NOR2X1 NOR2X1_370 ( .A(_3673_), .B(_3676_), .Y(_3677_) );
	NAND3X1 NAND3X1_155 ( .A(_3669_), .B(_3670_), .C(_3677_), .Y(_3678_) );
	AND2X2 AND2X2_68 ( .A(_3300_), .B(_3234_), .Y(_3679_) );
	AOI22X1 AOI22X1_499 ( .A(_3239_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_3679_), .Y(_3680_) );
	AND2X2 AND2X2_69 ( .A(_3298_), .B(_3263_), .Y(_3681_) );
	AND2X2 AND2X2_70 ( .A(_3306_), .B(_3263_), .Y(_3682_) );
	AOI22X1 AOI22X1_500 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_3682_), .C(_3681_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_3683_) );
	NAND2X1 NAND2X1_641 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_3391_), .Y(_3684_) );
	NAND2X1 NAND2X1_642 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_3364_), .Y(_3685_) );
	NAND2X1 NAND2X1_643 ( .A(_3684_), .B(_3685_), .Y(_3686_) );
	INVX1 INVX1_401 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_3687_) );
	NAND2X1 NAND2X1_644 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_3363_), .Y(_3688_) );
	OAI21X1 OAI21X1_106 ( .A(_3687_), .B(_3316_), .C(_3688_), .Y(_3689_) );
	NOR2X1 NOR2X1_371 ( .A(_3686_), .B(_3689_), .Y(_3690_) );
	NAND3X1 NAND3X1_156 ( .A(_3680_), .B(_3683_), .C(_3690_), .Y(_3691_) );
	NOR3X1 NOR3X1_266 ( .A(_3678_), .B(_3668_), .C(_3691_), .Y(_3692_) );
	INVX1 INVX1_402 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_3693_) );
	NAND2X1 NAND2X1_645 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_3279_), .Y(_3694_) );
	OAI21X1 OAI21X1_107 ( .A(_3284_), .B(_3693_), .C(_3694_), .Y(_3695_) );
	AOI21X1 AOI21X1_76 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_3259_), .C(_3695_), .Y(_3696_) );
	INVX1 INVX1_403 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_3697_) );
	INVX1 INVX1_404 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_3698_) );
	OAI22X1 OAI22X1_86 ( .A(_3603_), .B(_3698_), .C(_3697_), .D(_3254_), .Y(_3699_) );
	INVX1 INVX1_405 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_3700_) );
	NAND2X1 NAND2X1_646 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_3399_), .Y(_3701_) );
	OAI21X1 OAI21X1_108 ( .A(_3264_), .B(_3700_), .C(_3701_), .Y(_3702_) );
	NOR2X1 NOR2X1_372 ( .A(_3702_), .B(_3699_), .Y(_3703_) );
	INVX1 INVX1_406 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_3704_) );
	INVX1 INVX1_407 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_3705_) );
	OAI22X1 OAI22X1_87 ( .A(_3351_), .B(_3705_), .C(_3704_), .D(_3352_), .Y(_3706_) );
	INVX1 INVX1_408 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_3707_) );
	NAND2X1 NAND2X1_647 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_3398_), .Y(_3708_) );
	OAI21X1 OAI21X1_109 ( .A(_3707_), .B(_3334_), .C(_3708_), .Y(_3709_) );
	NOR2X1 NOR2X1_373 ( .A(_3709_), .B(_3706_), .Y(_3710_) );
	NAND3X1 NAND3X1_157 ( .A(_3696_), .B(_3710_), .C(_3703_), .Y(_3711_) );
	AOI22X1 AOI22X1_501 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_3356_), .C(_3357_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_3712_) );
	AOI22X1 AOI22X1_502 ( .A(_3359_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_3360_), .Y(_3713_) );
	NAND2X1 NAND2X1_648 ( .A(_3712_), .B(_3713_), .Y(_3714_) );
	AOI22X1 AOI22X1_503 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_3367_), .C(_3366_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_3715_) );
	AOI22X1 AOI22X1_504 ( .A(_3310_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_3317_), .Y(_3716_) );
	NAND2X1 NAND2X1_649 ( .A(_3715_), .B(_3716_), .Y(_3717_) );
	NOR2X1 NOR2X1_374 ( .A(_3714_), .B(_3717_), .Y(_3718_) );
	AOI22X1 AOI22X1_505 ( .A(_3371_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_3372_), .Y(_3719_) );
	AOI22X1 AOI22X1_506 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_3607_), .C(_3374_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_3720_) );
	NAND2X1 NAND2X1_650 ( .A(_3720_), .B(_3719_), .Y(_3721_) );
	AOI22X1 AOI22X1_507 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_3378_), .C(_3379_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_3722_) );
	AOI22X1 AOI22X1_508 ( .A(_3381_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_3382_), .Y(_3723_) );
	NAND2X1 NAND2X1_651 ( .A(_3723_), .B(_3722_), .Y(_3724_) );
	NOR2X1 NOR2X1_375 ( .A(_3721_), .B(_3724_), .Y(_3725_) );
	NAND2X1 NAND2X1_652 ( .A(_3725_), .B(_3718_), .Y(_3726_) );
	AOI22X1 AOI22X1_509 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_3388_), .C(_3289_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_3727_) );
	AOI22X1 AOI22X1_510 ( .A(_3312_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_3390_), .Y(_3728_) );
	NAND2X1 NAND2X1_653 ( .A(_3727_), .B(_3728_), .Y(_3729_) );
	AOI22X1 AOI22X1_511 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_3396_), .C(_3394_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_3730_) );
	AOI22X1 AOI22X1_512 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_3326_), .C(_3375_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_3731_) );
	NAND2X1 NAND2X1_654 ( .A(_3731_), .B(_3730_), .Y(_3732_) );
	NOR2X1 NOR2X1_376 ( .A(_3732_), .B(_3729_), .Y(_3733_) );
	AOI22X1 AOI22X1_513 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_3403_), .C(_3404_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_3734_) );
	NAND2X1 NAND2X1_655 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_3406_), .Y(_3735_) );
	NAND2X1 NAND2X1_656 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_3408_), .Y(_3736_) );
	NAND3X1 NAND3X1_158 ( .A(_3735_), .B(_3736_), .C(_3734_), .Y(_3737_) );
	AOI22X1 AOI22X1_514 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_3412_), .C(_3411_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_3738_) );
	AOI22X1 AOI22X1_515 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_3415_), .C(_3414_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_3739_) );
	NAND2X1 NAND2X1_657 ( .A(_3738_), .B(_3739_), .Y(_3740_) );
	NOR2X1 NOR2X1_377 ( .A(_3740_), .B(_3737_), .Y(_3741_) );
	NAND2X1 NAND2X1_658 ( .A(_3733_), .B(_3741_), .Y(_3742_) );
	NOR3X1 NOR3X1_267 ( .A(_3726_), .B(_3711_), .C(_3742_), .Y(_3743_) );
	NAND2X1 NAND2X1_659 ( .A(wData[59]), .B(_3445_), .Y(_3744_) );
	OAI21X1 OAI21X1_110 ( .A(_3229_), .B(wBusy_bF_buf4), .C(_3744_), .Y(_3745_) );
	NAND2X1 NAND2X1_660 ( .A(wData[7]), .B(_3436_), .Y(_3746_) );
	NAND2X1 NAND2X1_661 ( .A(wData[55]), .B(_3446_), .Y(_3747_) );
	AOI22X1 AOI22X1_516 ( .A(wData[63]), .B(_3448_), .C(_3438_), .D(wData[31]), .Y(_3748_) );
	NAND3X1 NAND3X1_159 ( .A(_3746_), .B(_3747_), .C(_3748_), .Y(_3749_) );
	OR2X2 OR2X2_36 ( .A(_3749_), .B(_3745_), .Y(_3750_) );
	INVX1 INVX1_409 ( .A(wData[51]), .Y(_3751_) );
	NAND2X1 NAND2X1_662 ( .A(wData[47]), .B(_3449_), .Y(_3752_) );
	OAI21X1 OAI21X1_111 ( .A(_3751_), .B(_3461_), .C(_3752_), .Y(_3753_) );
	AOI21X1 AOI21X1_77 ( .A(wData[3]), .B(_3456_), .C(_3753_), .Y(_3754_) );
	AOI22X1 AOI22X1_517 ( .A(_3462_), .B(wData[11]), .C(wData[15]), .D(_3463_), .Y(_3755_) );
	AOI22X1 AOI22X1_518 ( .A(_3425_), .B(wData[23]), .C(wData[27]), .D(_3432_), .Y(_3756_) );
	AND2X2 AND2X2_71 ( .A(_3755_), .B(_3756_), .Y(_3757_) );
	NAND2X1 NAND2X1_663 ( .A(wData[39]), .B(_3454_), .Y(_3758_) );
	NAND2X1 NAND2X1_664 ( .A(wData[43]), .B(_3452_), .Y(_3759_) );
	NAND2X1 NAND2X1_665 ( .A(_3758_), .B(_3759_), .Y(_3760_) );
	NAND2X1 NAND2X1_666 ( .A(wData[19]), .B(_3428_), .Y(_3761_) );
	NAND2X1 NAND2X1_667 ( .A(wData[35]), .B(_3442_), .Y(_3762_) );
	NAND2X1 NAND2X1_668 ( .A(_3761_), .B(_3762_), .Y(_3763_) );
	NOR2X1 NOR2X1_378 ( .A(_3760_), .B(_3763_), .Y(_3764_) );
	NAND3X1 NAND3X1_160 ( .A(_3757_), .B(_3754_), .C(_3764_), .Y(_3765_) );
	NOR2X1 NOR2X1_379 ( .A(_3750_), .B(_3765_), .Y(_3766_) );
	AOI21X1 AOI21X1_78 ( .A(_3692_), .B(_3743_), .C(_3766_), .Y(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_3_) );
	INVX1 INVX1_410 ( .A(wSelec[77]), .Y(_3767_) );
	NOR2X1 NOR2X1_380 ( .A(wBusy_bF_buf3), .B(_3767_), .Y(_3768_) );
	INVX1 INVX1_411 ( .A(_3768_), .Y(_3769_) );
	INVX1 INVX1_412 ( .A(wSelec[87]), .Y(_3770_) );
	NAND2X1 NAND2X1_669 ( .A(wSelec[86]), .B(_3770_), .Y(_3771_) );
	INVX2 INVX2_11 ( .A(_3771_), .Y(_3772_) );
	OR2X2 OR2X2_37 ( .A(wSelec[83]), .B(wSelec[82]), .Y(_3773_) );
	INVX1 INVX1_413 ( .A(wSelec[85]), .Y(_3774_) );
	NAND2X1 NAND2X1_670 ( .A(wSelec[84]), .B(_3774_), .Y(_3775_) );
	NOR2X1 NOR2X1_381 ( .A(_3773_), .B(_3775_), .Y(_3776_) );
	AND2X2 AND2X2_72 ( .A(_3776_), .B(_3772_), .Y(_3777_) );
	AOI21X1 AOI21X1_79 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_3777_), .C(_3769_), .Y(_3778_) );
	INVX1 INVX1_414 ( .A(wSelec[83]), .Y(_3779_) );
	NAND2X1 NAND2X1_671 ( .A(wSelec[82]), .B(_3779_), .Y(_3780_) );
	OR2X2 OR2X2_38 ( .A(wSelec[84]), .B(wSelec[85]), .Y(_3781_) );
	NOR2X1 NOR2X1_382 ( .A(_3781_), .B(_3780_), .Y(_3782_) );
	NAND2X1 NAND2X1_672 ( .A(_3772_), .B(_3782_), .Y(_3783_) );
	INVX1 INVX1_415 ( .A(_3783_), .Y(_3784_) );
	INVX1 INVX1_416 ( .A(wSelec[82]), .Y(_3785_) );
	NAND2X1 NAND2X1_673 ( .A(wSelec[83]), .B(_3785_), .Y(_3786_) );
	INVX1 INVX1_417 ( .A(wSelec[84]), .Y(_3787_) );
	NAND2X1 NAND2X1_674 ( .A(wSelec[85]), .B(_3787_), .Y(_3788_) );
	NOR2X1 NOR2X1_383 ( .A(_3786_), .B(_3788_), .Y(_3789_) );
	NAND2X1 NAND2X1_675 ( .A(wSelec[86]), .B(wSelec[87]), .Y(_3790_) );
	INVX1 INVX1_418 ( .A(_3790_), .Y(_3791_) );
	NAND2X1 NAND2X1_676 ( .A(_3791_), .B(_3789_), .Y(_3792_) );
	INVX1 INVX1_419 ( .A(_3792_), .Y(_3793_) );
	AOI22X1 AOI22X1_519 ( .A(_3784_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_3793_), .Y(_3794_) );
	OR2X2 OR2X2_39 ( .A(_3780_), .B(_3781_), .Y(_3795_) );
	OR2X2 OR2X2_40 ( .A(wSelec[86]), .B(wSelec[87]), .Y(_3796_) );
	NOR2X1 NOR2X1_384 ( .A(_3796_), .B(_3795_), .Y(_3797_) );
	NOR2X1 NOR2X1_385 ( .A(_3775_), .B(_3780_), .Y(_3798_) );
	INVX1 INVX1_420 ( .A(wSelec[86]), .Y(_3799_) );
	NAND2X1 NAND2X1_677 ( .A(wSelec[87]), .B(_3799_), .Y(_3800_) );
	INVX2 INVX2_12 ( .A(_3800_), .Y(_3801_) );
	NAND2X1 NAND2X1_678 ( .A(_3801_), .B(_3798_), .Y(_3802_) );
	INVX1 INVX1_421 ( .A(_3802_), .Y(_3803_) );
	AOI22X1 AOI22X1_520 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_3797_), .C(_3803_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_3804_) );
	NAND3X1 NAND3X1_161 ( .A(_3778_), .B(_3804_), .C(_3794_), .Y(_3805_) );
	NOR2X1 NOR2X1_386 ( .A(wSelec[83]), .B(wSelec[82]), .Y(_3806_) );
	NOR2X1 NOR2X1_387 ( .A(wSelec[84]), .B(wSelec[85]), .Y(_3807_) );
	NAND2X1 NAND2X1_679 ( .A(_3806_), .B(_3807_), .Y(_3808_) );
	NOR2X1 NOR2X1_388 ( .A(_3771_), .B(_3808_), .Y(_3809_) );
	NAND2X1 NAND2X1_680 ( .A(wSelec[83]), .B(wSelec[82]), .Y(_3810_) );
	NOR3X1 NOR3X1_268 ( .A(_3781_), .B(_3810_), .C(_3771_), .Y(_3811_) );
	AOI22X1 AOI22X1_521 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_3811_), .C(_3809_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_3812_) );
	INVX1 INVX1_422 ( .A(_3796_), .Y(_3813_) );
	NOR2X1 NOR2X1_389 ( .A(_3781_), .B(_3786_), .Y(_3814_) );
	AND2X2 AND2X2_73 ( .A(_3814_), .B(_3813_), .Y(_3815_) );
	NAND2X1 NAND2X1_681 ( .A(wSelec[84]), .B(wSelec[85]), .Y(_3816_) );
	NOR3X1 NOR3X1_269 ( .A(_3790_), .B(_3810_), .C(_3816_), .Y(_3817_) );
	AOI22X1 AOI22X1_522 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_3817_), .C(_3815_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_3818_) );
	INVX1 INVX1_423 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_3819_) );
	INVX1 INVX1_424 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_3820_) );
	NOR2X1 NOR2X1_390 ( .A(_3780_), .B(_3788_), .Y(_3821_) );
	NAND2X1 NAND2X1_682 ( .A(_3791_), .B(_3821_), .Y(_3822_) );
	NOR2X1 NOR2X1_391 ( .A(_3810_), .B(_3816_), .Y(_3823_) );
	NAND2X1 NAND2X1_683 ( .A(_3823_), .B(_3801_), .Y(_3824_) );
	OAI22X1 OAI22X1_88 ( .A(_3819_), .B(_3824_), .C(_3822_), .D(_3820_), .Y(_3825_) );
	INVX1 INVX1_425 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_3826_) );
	NOR3X1 NOR3X1_270 ( .A(_3771_), .B(_3786_), .C(_3788_), .Y(_3827_) );
	NAND2X1 NAND2X1_684 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_3827_), .Y(_3828_) );
	NOR2X1 NOR2X1_392 ( .A(_3810_), .B(_3775_), .Y(_3829_) );
	NAND2X1 NAND2X1_685 ( .A(_3801_), .B(_3829_), .Y(_3830_) );
	OAI21X1 OAI21X1_112 ( .A(_3826_), .B(_3830_), .C(_3828_), .Y(_3831_) );
	NOR2X1 NOR2X1_393 ( .A(_3825_), .B(_3831_), .Y(_3832_) );
	NAND3X1 NAND3X1_162 ( .A(_3812_), .B(_3818_), .C(_3832_), .Y(_3833_) );
	INVX1 INVX1_426 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_3834_) );
	INVX1 INVX1_427 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_3835_) );
	NOR2X1 NOR2X1_394 ( .A(_3775_), .B(_3786_), .Y(_3836_) );
	NAND2X1 NAND2X1_686 ( .A(_3772_), .B(_3836_), .Y(_3837_) );
	NOR2X1 NOR2X1_395 ( .A(_3773_), .B(_3788_), .Y(_3838_) );
	NAND2X1 NAND2X1_687 ( .A(_3772_), .B(_3838_), .Y(_3839_) );
	OAI22X1 OAI22X1_89 ( .A(_3839_), .B(_3834_), .C(_3835_), .D(_3837_), .Y(_3840_) );
	INVX1 INVX1_428 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_3841_) );
	INVX1 INVX1_429 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_3842_) );
	NAND2X1 NAND2X1_688 ( .A(_3801_), .B(_3836_), .Y(_3843_) );
	NOR2X1 NOR2X1_396 ( .A(_3810_), .B(_3781_), .Y(_3844_) );
	NAND2X1 NAND2X1_689 ( .A(_3801_), .B(_3844_), .Y(_3845_) );
	OAI22X1 OAI22X1_90 ( .A(_3841_), .B(_3845_), .C(_3843_), .D(_3842_), .Y(_3846_) );
	NOR2X1 NOR2X1_397 ( .A(_3846_), .B(_3840_), .Y(_3847_) );
	NOR3X1 NOR3X1_271 ( .A(_3780_), .B(_3816_), .C(_3800_), .Y(_3848_) );
	NAND2X1 NAND2X1_690 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_3848_), .Y(_3849_) );
	NOR3X1 NOR3X1_272 ( .A(_3788_), .B(_3810_), .C(_3800_), .Y(_3850_) );
	NAND2X1 NAND2X1_691 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_3850_), .Y(_3851_) );
	NAND2X1 NAND2X1_692 ( .A(_3849_), .B(_3851_), .Y(_3852_) );
	INVX1 INVX1_430 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_3853_) );
	NAND2X1 NAND2X1_693 ( .A(_3791_), .B(_3776_), .Y(_3854_) );
	NOR3X1 NOR3X1_273 ( .A(_3786_), .B(_3788_), .C(_3800_), .Y(_3855_) );
	NAND2X1 NAND2X1_694 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_3855_), .Y(_3856_) );
	OAI21X1 OAI21X1_113 ( .A(_3853_), .B(_3854_), .C(_3856_), .Y(_3857_) );
	NOR2X1 NOR2X1_398 ( .A(_3852_), .B(_3857_), .Y(_3858_) );
	NAND2X1 NAND2X1_695 ( .A(_3847_), .B(_3858_), .Y(_3859_) );
	NOR3X1 NOR3X1_274 ( .A(_3805_), .B(_3859_), .C(_3833_), .Y(_3860_) );
	NAND2X1 NAND2X1_696 ( .A(_3772_), .B(_3829_), .Y(_3861_) );
	INVX1 INVX1_431 ( .A(_3861_), .Y(_3862_) );
	INVX1 INVX1_432 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_3863_) );
	NOR3X1 NOR3X1_275 ( .A(_3773_), .B(_3796_), .C(_3775_), .Y(_3864_) );
	NAND2X1 NAND2X1_697 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_3864_), .Y(_3865_) );
	NAND2X1 NAND2X1_698 ( .A(_3813_), .B(_3836_), .Y(_3866_) );
	OAI21X1 OAI21X1_114 ( .A(_3866_), .B(_3863_), .C(_3865_), .Y(_3867_) );
	AOI21X1 AOI21X1_80 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_3862_), .C(_3867_), .Y(_3868_) );
	INVX1 INVX1_433 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_3869_) );
	INVX1 INVX1_434 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_3870_) );
	NOR2X1 NOR2X1_399 ( .A(_3816_), .B(_3773_), .Y(_3871_) );
	NAND2X1 NAND2X1_699 ( .A(_3772_), .B(_3871_), .Y(_3872_) );
	NAND2X1 NAND2X1_700 ( .A(_3813_), .B(_3798_), .Y(_3873_) );
	OAI22X1 OAI22X1_91 ( .A(_3870_), .B(_3872_), .C(_3873_), .D(_3869_), .Y(_3874_) );
	INVX1 INVX1_435 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_3875_) );
	INVX1 INVX1_436 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_3876_) );
	NAND2X1 NAND2X1_701 ( .A(_3772_), .B(_3798_), .Y(_3877_) );
	NAND2X1 NAND2X1_702 ( .A(_3813_), .B(_3844_), .Y(_3878_) );
	OAI22X1 OAI22X1_92 ( .A(_3875_), .B(_3878_), .C(_3877_), .D(_3876_), .Y(_3879_) );
	NOR2X1 NOR2X1_400 ( .A(_3874_), .B(_3879_), .Y(_3880_) );
	INVX1 INVX1_437 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_3881_) );
	NOR3X1 NOR3X1_276 ( .A(_3796_), .B(_3810_), .C(_3775_), .Y(_3882_) );
	NAND2X1 NAND2X1_703 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_3882_), .Y(_3883_) );
	OR2X2 OR2X2_41 ( .A(_3808_), .B(_3790_), .Y(_3884_) );
	OAI21X1 OAI21X1_115 ( .A(_3881_), .B(_3884_), .C(_3883_), .Y(_3885_) );
	INVX1 INVX1_438 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_3886_) );
	INVX1 INVX1_439 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_3887_) );
	NOR2X1 NOR2X1_401 ( .A(_3816_), .B(_3786_), .Y(_3888_) );
	NAND2X1 NAND2X1_704 ( .A(_3772_), .B(_3888_), .Y(_3889_) );
	NAND2X1 NAND2X1_705 ( .A(_3791_), .B(_3782_), .Y(_3890_) );
	OAI22X1 OAI22X1_93 ( .A(_3889_), .B(_3887_), .C(_3886_), .D(_3890_), .Y(_3891_) );
	NOR2X1 NOR2X1_402 ( .A(_3885_), .B(_3891_), .Y(_3892_) );
	NAND3X1 NAND3X1_163 ( .A(_3868_), .B(_3892_), .C(_3880_), .Y(_3893_) );
	NOR3X1 NOR3X1_277 ( .A(_3773_), .B(_3781_), .C(_3796_), .Y(_3894_) );
	NOR3X1 NOR3X1_278 ( .A(_3790_), .B(_3816_), .C(_3780_), .Y(_3895_) );
	AOI22X1 AOI22X1_523 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_3894_), .C(_3895_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_3896_) );
	NOR3X1 NOR3X1_279 ( .A(_3790_), .B(_3816_), .C(_3786_), .Y(_3897_) );
	NOR3X1 NOR3X1_280 ( .A(_3790_), .B(_3810_), .C(_3788_), .Y(_3898_) );
	AOI22X1 AOI22X1_524 ( .A(_3897_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_3898_), .Y(_3899_) );
	NAND2X1 NAND2X1_706 ( .A(_3896_), .B(_3899_), .Y(_3900_) );
	NOR3X1 NOR3X1_281 ( .A(_3788_), .B(_3773_), .C(_3800_), .Y(_3901_) );
	NOR3X1 NOR3X1_282 ( .A(_3780_), .B(_3788_), .C(_3800_), .Y(_3902_) );
	AOI22X1 AOI22X1_525 ( .A(_3901_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_3902_), .Y(_3903_) );
	NOR3X1 NOR3X1_283 ( .A(_3771_), .B(_3816_), .C(_3780_), .Y(_3904_) );
	NOR3X1 NOR3X1_284 ( .A(_3810_), .B(_3816_), .C(_3771_), .Y(_3905_) );
	AOI22X1 AOI22X1_526 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_3905_), .C(_3904_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_3906_) );
	NAND2X1 NAND2X1_707 ( .A(_3906_), .B(_3903_), .Y(_3907_) );
	NOR2X1 NOR2X1_403 ( .A(_3900_), .B(_3907_), .Y(_3908_) );
	NOR3X1 NOR3X1_285 ( .A(_3796_), .B(_3816_), .C(_3780_), .Y(_3909_) );
	NOR3X1 NOR3X1_286 ( .A(_3796_), .B(_3816_), .C(_3786_), .Y(_3910_) );
	AOI22X1 AOI22X1_527 ( .A(_3909_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_3910_), .Y(_3911_) );
	NOR3X1 NOR3X1_287 ( .A(_3796_), .B(_3810_), .C(_3788_), .Y(_3912_) );
	NOR3X1 NOR3X1_288 ( .A(_3771_), .B(_3781_), .C(_3786_), .Y(_3913_) );
	AOI22X1 AOI22X1_528 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_3912_), .C(_3913_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_3914_) );
	NAND2X1 NAND2X1_708 ( .A(_3911_), .B(_3914_), .Y(_3915_) );
	NOR3X1 NOR3X1_289 ( .A(_3810_), .B(_3816_), .C(_3796_), .Y(_3916_) );
	NOR3X1 NOR3X1_290 ( .A(_3786_), .B(_3781_), .C(_3800_), .Y(_3917_) );
	AOI22X1 AOI22X1_529 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_3916_), .C(_3917_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_3918_) );
	NOR3X1 NOR3X1_291 ( .A(_3773_), .B(_3781_), .C(_3800_), .Y(_3919_) );
	NOR3X1 NOR3X1_292 ( .A(_3773_), .B(_3816_), .C(_3800_), .Y(_3920_) );
	AOI22X1 AOI22X1_530 ( .A(_3919_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_3920_), .Y(_3921_) );
	NAND2X1 NAND2X1_709 ( .A(_3921_), .B(_3918_), .Y(_3922_) );
	NOR2X1 NOR2X1_404 ( .A(_3915_), .B(_3922_), .Y(_3923_) );
	NAND2X1 NAND2X1_710 ( .A(_3923_), .B(_3908_), .Y(_3924_) );
	NOR3X1 NOR3X1_293 ( .A(_3771_), .B(_3810_), .C(_3788_), .Y(_3925_) );
	NOR3X1 NOR3X1_294 ( .A(_3781_), .B(_3790_), .C(_3786_), .Y(_3926_) );
	AOI22X1 AOI22X1_531 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_3926_), .C(_3925_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_3927_) );
	NOR3X1 NOR3X1_295 ( .A(_3775_), .B(_3773_), .C(_3800_), .Y(_3928_) );
	NOR3X1 NOR3X1_296 ( .A(_3786_), .B(_3816_), .C(_3800_), .Y(_3929_) );
	AOI22X1 AOI22X1_532 ( .A(_3928_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_3929_), .Y(_3930_) );
	NAND2X1 NAND2X1_711 ( .A(_3927_), .B(_3930_), .Y(_3931_) );
	NOR3X1 NOR3X1_297 ( .A(_3771_), .B(_3780_), .C(_3788_), .Y(_3932_) );
	NAND2X1 NAND2X1_712 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_3932_), .Y(_3933_) );
	NOR3X1 NOR3X1_298 ( .A(_3790_), .B(_3810_), .C(_3775_), .Y(_3934_) );
	NAND2X1 NAND2X1_713 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_3934_), .Y(_3935_) );
	NOR3X1 NOR3X1_299 ( .A(_3773_), .B(_3816_), .C(_3796_), .Y(_3936_) );
	NOR3X1 NOR3X1_300 ( .A(_3773_), .B(_3790_), .C(_3788_), .Y(_3937_) );
	AOI22X1 AOI22X1_533 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_3936_), .C(_3937_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_3938_) );
	NAND3X1 NAND3X1_164 ( .A(_3933_), .B(_3935_), .C(_3938_), .Y(_3939_) );
	NOR2X1 NOR2X1_405 ( .A(_3939_), .B(_3931_), .Y(_3940_) );
	NOR3X1 NOR3X1_301 ( .A(_3773_), .B(_3796_), .C(_3788_), .Y(_3941_) );
	NOR3X1 NOR3X1_302 ( .A(_3775_), .B(_3790_), .C(_3780_), .Y(_3942_) );
	AOI22X1 AOI22X1_534 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_3941_), .C(_3942_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_3943_) );
	NOR3X1 NOR3X1_303 ( .A(_3775_), .B(_3790_), .C(_3786_), .Y(_3944_) );
	NAND2X1 NAND2X1_714 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_3944_), .Y(_3945_) );
	NOR3X1 NOR3X1_304 ( .A(_3780_), .B(_3781_), .C(_3800_), .Y(_3946_) );
	NAND2X1 NAND2X1_715 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_3946_), .Y(_3947_) );
	NAND3X1 NAND3X1_165 ( .A(_3945_), .B(_3947_), .C(_3943_), .Y(_3948_) );
	NOR3X1 NOR3X1_305 ( .A(_3780_), .B(_3796_), .C(_3788_), .Y(_3949_) );
	NOR3X1 NOR3X1_306 ( .A(_3790_), .B(_3816_), .C(_3773_), .Y(_3950_) );
	AOI22X1 AOI22X1_535 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_3950_), .C(_3949_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_3951_) );
	NOR3X1 NOR3X1_307 ( .A(_3786_), .B(_3796_), .C(_3788_), .Y(_3952_) );
	NOR3X1 NOR3X1_308 ( .A(_3790_), .B(_3810_), .C(_3781_), .Y(_3953_) );
	AOI22X1 AOI22X1_536 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_3953_), .C(_3952_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_3954_) );
	NAND2X1 NAND2X1_716 ( .A(_3951_), .B(_3954_), .Y(_3955_) );
	NOR2X1 NOR2X1_406 ( .A(_3955_), .B(_3948_), .Y(_3956_) );
	NAND2X1 NAND2X1_717 ( .A(_3940_), .B(_3956_), .Y(_3957_) );
	NOR3X1 NOR3X1_309 ( .A(_3924_), .B(_3893_), .C(_3957_), .Y(_3958_) );
	INVX1 INVX1_440 ( .A(wSelec[79]), .Y(_3959_) );
	NAND2X1 NAND2X1_718 ( .A(wSelec[78]), .B(_3959_), .Y(_3960_) );
	INVX1 INVX1_441 ( .A(wSelec[81]), .Y(_3961_) );
	NAND2X1 NAND2X1_719 ( .A(wSelec[80]), .B(_3961_), .Y(_3962_) );
	NOR2X1 NOR2X1_407 ( .A(_3960_), .B(_3962_), .Y(_3963_) );
	NOR2X1 NOR2X1_408 ( .A(wSelec[79]), .B(wSelec[78]), .Y(_3964_) );
	INVX1 INVX1_442 ( .A(_3964_), .Y(_3965_) );
	NOR2X1 NOR2X1_409 ( .A(_3962_), .B(_3965_), .Y(_3966_) );
	AOI22X1 AOI22X1_537 ( .A(wData[20]), .B(_3963_), .C(_3966_), .D(wData[16]), .Y(_3967_) );
	INVX1 INVX1_443 ( .A(wSelec[78]), .Y(_3968_) );
	NAND2X1 NAND2X1_720 ( .A(wSelec[79]), .B(_3968_), .Y(_3969_) );
	NOR2X1 NOR2X1_410 ( .A(_3969_), .B(_3962_), .Y(_3970_) );
	NAND2X1 NAND2X1_721 ( .A(wData[24]), .B(_3970_), .Y(_3971_) );
	INVX1 INVX1_444 ( .A(wSelec[80]), .Y(_3972_) );
	NAND2X1 NAND2X1_722 ( .A(_3972_), .B(_3961_), .Y(_3973_) );
	NOR2X1 NOR2X1_411 ( .A(_3960_), .B(_3973_), .Y(_3974_) );
	NAND2X1 NAND2X1_723 ( .A(wSelec[79]), .B(wSelec[78]), .Y(_3975_) );
	NOR2X1 NOR2X1_412 ( .A(_3975_), .B(_3962_), .Y(_3976_) );
	AOI22X1 AOI22X1_538 ( .A(_3976_), .B(wData[28]), .C(wData[4]), .D(_3974_), .Y(_3977_) );
	NAND3X1 NAND3X1_166 ( .A(_3971_), .B(_3977_), .C(_3967_), .Y(_3978_) );
	NAND2X1 NAND2X1_724 ( .A(wSelec[81]), .B(_3972_), .Y(_3979_) );
	NOR2X1 NOR2X1_413 ( .A(_3979_), .B(_3965_), .Y(_3980_) );
	NAND2X1 NAND2X1_725 ( .A(wData[32]), .B(_3980_), .Y(_3981_) );
	NAND2X1 NAND2X1_726 ( .A(wSelec[80]), .B(wSelec[81]), .Y(_3982_) );
	NOR2X1 NOR2X1_414 ( .A(_3982_), .B(_3969_), .Y(_3983_) );
	NOR2X1 NOR2X1_415 ( .A(_3982_), .B(_3960_), .Y(_3984_) );
	AOI22X1 AOI22X1_539 ( .A(_3983_), .B(wData[56]), .C(wData[52]), .D(_3984_), .Y(_3985_) );
	NOR2X1 NOR2X1_416 ( .A(_3975_), .B(_3982_), .Y(_3986_) );
	NOR2X1 NOR2X1_417 ( .A(_3975_), .B(_3979_), .Y(_3987_) );
	AOI22X1 AOI22X1_540 ( .A(wData[60]), .B(_3986_), .C(_3987_), .D(wData[44]), .Y(_3988_) );
	NAND3X1 NAND3X1_167 ( .A(_3981_), .B(_3988_), .C(_3985_), .Y(_3989_) );
	NOR2X1 NOR2X1_418 ( .A(_3969_), .B(_3979_), .Y(_3990_) );
	NAND2X1 NAND2X1_727 ( .A(wData[40]), .B(_3990_), .Y(_3991_) );
	NOR2X1 NOR2X1_419 ( .A(_3979_), .B(_3960_), .Y(_3992_) );
	NAND2X1 NAND2X1_728 ( .A(wData[36]), .B(_3992_), .Y(_3993_) );
	NOR2X1 NOR2X1_420 ( .A(_3973_), .B(_3965_), .Y(_3994_) );
	NAND2X1 NAND2X1_729 ( .A(wData[0]), .B(_3994_), .Y(_3995_) );
	NAND3X1 NAND3X1_168 ( .A(_3991_), .B(_3993_), .C(_3995_), .Y(_3996_) );
	INVX1 INVX1_445 ( .A(wData[48]), .Y(_3997_) );
	NOR2X1 NOR2X1_421 ( .A(_3972_), .B(_3961_), .Y(_3998_) );
	NAND2X1 NAND2X1_730 ( .A(_3964_), .B(_3998_), .Y(_3999_) );
	NOR2X1 NOR2X1_422 ( .A(_3969_), .B(_3973_), .Y(_4000_) );
	NOR2X1 NOR2X1_423 ( .A(_3975_), .B(_3973_), .Y(_4001_) );
	AOI22X1 AOI22X1_541 ( .A(_4000_), .B(wData[8]), .C(wData[12]), .D(_4001_), .Y(_4002_) );
	OAI21X1 OAI21X1_116 ( .A(_3997_), .B(_3999_), .C(_4002_), .Y(_4003_) );
	OR2X2 OR2X2_42 ( .A(_4003_), .B(_3996_), .Y(_4004_) );
	NOR3X1 NOR3X1_310 ( .A(_3978_), .B(_3989_), .C(_4004_), .Y(_4005_) );
	AND2X2 AND2X2_74 ( .A(_4005_), .B(_3769_), .Y(_4006_) );
	AOI21X1 AOI21X1_81 ( .A(_3860_), .B(_3958_), .C(_4006_), .Y(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_0_) );
	INVX1 INVX1_446 ( .A(_3877_), .Y(_4007_) );
	AOI21X1 AOI21X1_82 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_4007_), .C(_3769_), .Y(_4008_) );
	AOI22X1 AOI22X1_542 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_3777_), .C(_3793_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_4009_) );
	AOI22X1 AOI22X1_543 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_3797_), .C(_3803_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_4010_) );
	NAND3X1 NAND3X1_169 ( .A(_4008_), .B(_4009_), .C(_4010_), .Y(_4011_) );
	INVX1 INVX1_447 ( .A(_3837_), .Y(_4012_) );
	AOI22X1 AOI22X1_544 ( .A(_3862_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_4012_), .Y(_4013_) );
	AOI22X1 AOI22X1_545 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_3936_), .C(_3815_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_4014_) );
	INVX1 INVX1_448 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_4015_) );
	INVX1 INVX1_449 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_4016_) );
	OAI22X1 OAI22X1_94 ( .A(_4015_), .B(_3824_), .C(_3822_), .D(_4016_), .Y(_4017_) );
	INVX1 INVX1_450 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_4018_) );
	NAND2X1 NAND2X1_731 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_3925_), .Y(_4019_) );
	OAI21X1 OAI21X1_117 ( .A(_4018_), .B(_3830_), .C(_4019_), .Y(_4020_) );
	NOR2X1 NOR2X1_424 ( .A(_4017_), .B(_4020_), .Y(_4021_) );
	NAND3X1 NAND3X1_170 ( .A(_4013_), .B(_4014_), .C(_4021_), .Y(_4022_) );
	INVX1 INVX1_451 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_4023_) );
	NAND2X1 NAND2X1_732 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_3809_), .Y(_4024_) );
	OAI21X1 OAI21X1_118 ( .A(_4023_), .B(_3839_), .C(_4024_), .Y(_4025_) );
	INVX1 INVX1_452 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_4026_) );
	INVX1 INVX1_453 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_4027_) );
	OAI22X1 OAI22X1_95 ( .A(_4026_), .B(_3845_), .C(_3843_), .D(_4027_), .Y(_4028_) );
	NOR2X1 NOR2X1_425 ( .A(_4028_), .B(_4025_), .Y(_4029_) );
	AOI22X1 AOI22X1_546 ( .A(_3929_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_3902_), .Y(_4030_) );
	AND2X2 AND2X2_75 ( .A(_3776_), .B(_3791_), .Y(_4031_) );
	AOI22X1 AOI22X1_547 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_3901_), .C(_4031_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_4032_) );
	NAND3X1 NAND3X1_171 ( .A(_4030_), .B(_4032_), .C(_4029_), .Y(_4033_) );
	NOR3X1 NOR3X1_311 ( .A(_4033_), .B(_4011_), .C(_4022_), .Y(_4034_) );
	INVX1 INVX1_454 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_4035_) );
	NAND2X1 NAND2X1_733 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_3864_), .Y(_4036_) );
	OAI21X1 OAI21X1_119 ( .A(_3866_), .B(_4035_), .C(_4036_), .Y(_4037_) );
	AOI21X1 AOI21X1_83 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_3913_), .C(_4037_), .Y(_4038_) );
	INVX1 INVX1_455 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_4039_) );
	INVX1 INVX1_456 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_4040_) );
	OAI22X1 OAI22X1_96 ( .A(_4040_), .B(_3872_), .C(_3873_), .D(_4039_), .Y(_4041_) );
	INVX1 INVX1_457 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_4042_) );
	NAND2X1 NAND2X1_734 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_3882_), .Y(_4043_) );
	OAI21X1 OAI21X1_120 ( .A(_3783_), .B(_4042_), .C(_4043_), .Y(_4044_) );
	NOR2X1 NOR2X1_426 ( .A(_4044_), .B(_4041_), .Y(_4045_) );
	INVX1 INVX1_458 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_4046_) );
	INVX1 INVX1_459 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_4047_) );
	OAI22X1 OAI22X1_97 ( .A(_3878_), .B(_4047_), .C(_3884_), .D(_4046_), .Y(_4048_) );
	INVX1 INVX1_460 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_4049_) );
	NOR2X1 NOR2X1_427 ( .A(_4049_), .B(_3889_), .Y(_4050_) );
	INVX1 INVX1_461 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_4051_) );
	NOR2X1 NOR2X1_428 ( .A(_4051_), .B(_3890_), .Y(_4052_) );
	NOR3X1 NOR3X1_312 ( .A(_4050_), .B(_4048_), .C(_4052_), .Y(_4053_) );
	NAND3X1 NAND3X1_172 ( .A(_4045_), .B(_4038_), .C(_4053_), .Y(_4054_) );
	AOI22X1 AOI22X1_548 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_3894_), .C(_3895_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_4055_) );
	AOI22X1 AOI22X1_549 ( .A(_3897_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_3898_), .Y(_4056_) );
	NAND2X1 NAND2X1_735 ( .A(_4055_), .B(_4056_), .Y(_4057_) );
	AOI22X1 AOI22X1_550 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_3905_), .C(_3904_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_4058_) );
	AOI22X1 AOI22X1_551 ( .A(_3848_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_3855_), .Y(_4059_) );
	NAND2X1 NAND2X1_736 ( .A(_4058_), .B(_4059_), .Y(_4060_) );
	NOR2X1 NOR2X1_429 ( .A(_4057_), .B(_4060_), .Y(_4061_) );
	AOI22X1 AOI22X1_552 ( .A(_3909_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_3910_), .Y(_4062_) );
	AOI22X1 AOI22X1_553 ( .A(_3811_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_3912_), .Y(_4063_) );
	NAND2X1 NAND2X1_737 ( .A(_4062_), .B(_4063_), .Y(_4064_) );
	AOI22X1 AOI22X1_554 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_3916_), .C(_3917_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_4065_) );
	AOI22X1 AOI22X1_555 ( .A(_3919_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_3920_), .Y(_4066_) );
	NAND2X1 NAND2X1_738 ( .A(_4066_), .B(_4065_), .Y(_4067_) );
	NOR2X1 NOR2X1_430 ( .A(_4064_), .B(_4067_), .Y(_4068_) );
	NAND2X1 NAND2X1_739 ( .A(_4068_), .B(_4061_), .Y(_4069_) );
	AOI22X1 AOI22X1_556 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_3926_), .C(_3827_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_4070_) );
	AOI22X1 AOI22X1_557 ( .A(_3850_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_3928_), .Y(_4071_) );
	NAND2X1 NAND2X1_740 ( .A(_4070_), .B(_4071_), .Y(_4072_) );
	AOI22X1 AOI22X1_558 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_3817_), .C(_3937_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_4073_) );
	NAND2X1 NAND2X1_741 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_3932_), .Y(_4074_) );
	NAND2X1 NAND2X1_742 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_3934_), .Y(_4075_) );
	NAND3X1 NAND3X1_173 ( .A(_4074_), .B(_4075_), .C(_4073_), .Y(_4076_) );
	NOR2X1 NOR2X1_431 ( .A(_4076_), .B(_4072_), .Y(_4077_) );
	AOI22X1 AOI22X1_559 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_3941_), .C(_3942_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_4078_) );
	NAND2X1 NAND2X1_743 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_3944_), .Y(_4079_) );
	NAND2X1 NAND2X1_744 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_3946_), .Y(_4080_) );
	NAND3X1 NAND3X1_174 ( .A(_4079_), .B(_4080_), .C(_4078_), .Y(_4081_) );
	AOI22X1 AOI22X1_560 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_3950_), .C(_3949_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_4082_) );
	AOI22X1 AOI22X1_561 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_3953_), .C(_3952_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_4083_) );
	NAND2X1 NAND2X1_745 ( .A(_4082_), .B(_4083_), .Y(_4084_) );
	NOR2X1 NOR2X1_432 ( .A(_4084_), .B(_4081_), .Y(_4085_) );
	NAND2X1 NAND2X1_746 ( .A(_4077_), .B(_4085_), .Y(_4086_) );
	NOR3X1 NOR3X1_313 ( .A(_4069_), .B(_4054_), .C(_4086_), .Y(_4087_) );
	AOI21X1 AOI21X1_84 ( .A(wData[21]), .B(_3963_), .C(_3768_), .Y(_4088_) );
	AOI22X1 AOI22X1_562 ( .A(_3966_), .B(wData[17]), .C(wData[1]), .D(_3994_), .Y(_4089_) );
	AOI22X1 AOI22X1_563 ( .A(_3987_), .B(wData[45]), .C(wData[25]), .D(_3970_), .Y(_4090_) );
	NAND3X1 NAND3X1_175 ( .A(_4088_), .B(_4090_), .C(_4089_), .Y(_4091_) );
	NAND3X1 NAND3X1_176 ( .A(wData[49]), .B(_3964_), .C(_3998_), .Y(_4092_) );
	AOI22X1 AOI22X1_564 ( .A(wData[61]), .B(_3986_), .C(_3974_), .D(wData[5]), .Y(_4093_) );
	AND2X2 AND2X2_76 ( .A(_4093_), .B(_4092_), .Y(_4094_) );
	AOI22X1 AOI22X1_565 ( .A(_3983_), .B(wData[57]), .C(wData[41]), .D(_3990_), .Y(_4095_) );
	AOI22X1 AOI22X1_566 ( .A(wData[53]), .B(_3984_), .C(_3980_), .D(wData[33]), .Y(_4096_) );
	AND2X2 AND2X2_77 ( .A(_4096_), .B(_4095_), .Y(_4097_) );
	AOI22X1 AOI22X1_567 ( .A(_4000_), .B(wData[9]), .C(wData[13]), .D(_4001_), .Y(_4098_) );
	AOI22X1 AOI22X1_568 ( .A(_3976_), .B(wData[29]), .C(wData[37]), .D(_3992_), .Y(_4099_) );
	AND2X2 AND2X2_78 ( .A(_4098_), .B(_4099_), .Y(_4100_) );
	NAND3X1 NAND3X1_177 ( .A(_4094_), .B(_4100_), .C(_4097_), .Y(_4101_) );
	NOR2X1 NOR2X1_433 ( .A(_4091_), .B(_4101_), .Y(_4102_) );
	AOI21X1 AOI21X1_85 ( .A(_4034_), .B(_4087_), .C(_4102_), .Y(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_1_) );
	AOI21X1 AOI21X1_86 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_4007_), .C(_3769_), .Y(_4103_) );
	INVX1 INVX1_462 ( .A(_3866_), .Y(_4104_) );
	AOI22X1 AOI22X1_569 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_3777_), .C(_4104_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_4105_) );
	INVX1 INVX1_463 ( .A(_3878_), .Y(_4106_) );
	AOI22X1 AOI22X1_570 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_3913_), .C(_4106_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_4107_) );
	NAND3X1 NAND3X1_178 ( .A(_4107_), .B(_4103_), .C(_4105_), .Y(_4108_) );
	AOI22X1 AOI22X1_571 ( .A(_3862_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_4012_), .Y(_4109_) );
	AOI22X1 AOI22X1_572 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_3811_), .C(_3784_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_4110_) );
	INVX1 INVX1_464 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_4111_) );
	NAND2X1 NAND2X1_747 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_3901_), .Y(_4112_) );
	OAI21X1 OAI21X1_121 ( .A(_4111_), .B(_3873_), .C(_4112_), .Y(_4113_) );
	INVX1 INVX1_465 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_4114_) );
	NAND2X1 NAND2X1_748 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_3827_), .Y(_4115_) );
	OAI21X1 OAI21X1_122 ( .A(_4114_), .B(_3830_), .C(_4115_), .Y(_4116_) );
	NOR2X1 NOR2X1_434 ( .A(_4113_), .B(_4116_), .Y(_4117_) );
	NAND3X1 NAND3X1_179 ( .A(_4109_), .B(_4110_), .C(_4117_), .Y(_4118_) );
	INVX1 INVX1_466 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_4119_) );
	NAND2X1 NAND2X1_749 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_3809_), .Y(_4120_) );
	OAI21X1 OAI21X1_123 ( .A(_4119_), .B(_3839_), .C(_4120_), .Y(_4121_) );
	INVX1 INVX1_467 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_4122_) );
	INVX1 INVX1_468 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_4123_) );
	OAI22X1 OAI22X1_98 ( .A(_4122_), .B(_3845_), .C(_3843_), .D(_4123_), .Y(_4124_) );
	NOR2X1 NOR2X1_435 ( .A(_4124_), .B(_4121_), .Y(_4125_) );
	AOI22X1 AOI22X1_573 ( .A(_3929_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_3902_), .Y(_4126_) );
	AND2X2 AND2X2_79 ( .A(_3801_), .B(_3823_), .Y(_4127_) );
	AOI22X1 AOI22X1_574 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_4127_), .C(_4031_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_4128_) );
	NAND3X1 NAND3X1_180 ( .A(_4126_), .B(_4128_), .C(_4125_), .Y(_4129_) );
	NOR3X1 NOR3X1_314 ( .A(_4129_), .B(_4108_), .C(_4118_), .Y(_4130_) );
	INVX1 INVX1_469 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_4131_) );
	NOR3X1 NOR3X1_315 ( .A(_4131_), .B(_3796_), .C(_3795_), .Y(_4132_) );
	AND2X2 AND2X2_80 ( .A(_3817_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_4133_) );
	AND2X2 AND2X2_81 ( .A(_3937_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_4134_) );
	NOR3X1 NOR3X1_316 ( .A(_4134_), .B(_4133_), .C(_4132_), .Y(_4135_) );
	INVX1 INVX1_470 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_4136_) );
	INVX1 INVX1_471 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_4137_) );
	OAI22X1 OAI22X1_99 ( .A(_4137_), .B(_3872_), .C(_3822_), .D(_4136_), .Y(_4138_) );
	INVX1 INVX1_472 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_4139_) );
	INVX1 INVX1_473 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_4140_) );
	NAND2X1 NAND2X1_750 ( .A(_3813_), .B(_3814_), .Y(_4141_) );
	OAI22X1 OAI22X1_100 ( .A(_4141_), .B(_4140_), .C(_4139_), .D(_3792_), .Y(_4142_) );
	NOR2X1 NOR2X1_436 ( .A(_4138_), .B(_4142_), .Y(_4143_) );
	INVX1 INVX1_474 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_4144_) );
	NOR3X1 NOR3X1_317 ( .A(_3773_), .B(_3790_), .C(_3781_), .Y(_4145_) );
	NAND2X1 NAND2X1_751 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_4145_), .Y(_4146_) );
	OAI21X1 OAI21X1_124 ( .A(_3802_), .B(_4144_), .C(_4146_), .Y(_4147_) );
	INVX1 INVX1_475 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_4148_) );
	INVX1 INVX1_476 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_4149_) );
	OAI22X1 OAI22X1_101 ( .A(_3889_), .B(_4149_), .C(_4148_), .D(_3890_), .Y(_4150_) );
	NOR2X1 NOR2X1_437 ( .A(_4147_), .B(_4150_), .Y(_4151_) );
	NAND3X1 NAND3X1_181 ( .A(_4135_), .B(_4151_), .C(_4143_), .Y(_4152_) );
	AOI22X1 AOI22X1_575 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_3894_), .C(_3895_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_4153_) );
	AOI22X1 AOI22X1_576 ( .A(_3897_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_3898_), .Y(_4154_) );
	NAND2X1 NAND2X1_752 ( .A(_4153_), .B(_4154_), .Y(_4155_) );
	AOI22X1 AOI22X1_577 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_3905_), .C(_3904_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_4156_) );
	AOI22X1 AOI22X1_578 ( .A(_3848_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_3855_), .Y(_4157_) );
	NAND2X1 NAND2X1_753 ( .A(_4156_), .B(_4157_), .Y(_4158_) );
	NOR2X1 NOR2X1_438 ( .A(_4155_), .B(_4158_), .Y(_4159_) );
	AOI22X1 AOI22X1_579 ( .A(_3909_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_3910_), .Y(_4160_) );
	AOI22X1 AOI22X1_580 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_3936_), .C(_3912_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_4161_) );
	NAND2X1 NAND2X1_754 ( .A(_4161_), .B(_4160_), .Y(_4162_) );
	AOI22X1 AOI22X1_581 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_3916_), .C(_3917_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_4163_) );
	AOI22X1 AOI22X1_582 ( .A(_3919_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_3920_), .Y(_4164_) );
	NAND2X1 NAND2X1_755 ( .A(_4164_), .B(_4163_), .Y(_4165_) );
	NOR2X1 NOR2X1_439 ( .A(_4162_), .B(_4165_), .Y(_4166_) );
	NAND2X1 NAND2X1_756 ( .A(_4166_), .B(_4159_), .Y(_4167_) );
	AOI22X1 AOI22X1_583 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_3926_), .C(_3925_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_4168_) );
	AOI22X1 AOI22X1_584 ( .A(_3850_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_3928_), .Y(_4169_) );
	NAND2X1 NAND2X1_757 ( .A(_4168_), .B(_4169_), .Y(_4170_) );
	AOI22X1 AOI22X1_585 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_3934_), .C(_3932_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_4171_) );
	AOI22X1 AOI22X1_586 ( .A(_3864_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_3882_), .Y(_4172_) );
	NAND2X1 NAND2X1_758 ( .A(_4172_), .B(_4171_), .Y(_4173_) );
	NOR2X1 NOR2X1_440 ( .A(_4173_), .B(_4170_), .Y(_4174_) );
	AOI22X1 AOI22X1_587 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_3941_), .C(_3942_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_4175_) );
	NAND2X1 NAND2X1_759 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_3944_), .Y(_4176_) );
	NAND2X1 NAND2X1_760 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_3946_), .Y(_4177_) );
	NAND3X1 NAND3X1_182 ( .A(_4176_), .B(_4177_), .C(_4175_), .Y(_4178_) );
	AOI22X1 AOI22X1_588 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_3950_), .C(_3949_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_4179_) );
	AOI22X1 AOI22X1_589 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_3953_), .C(_3952_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_4180_) );
	NAND2X1 NAND2X1_761 ( .A(_4179_), .B(_4180_), .Y(_4181_) );
	NOR2X1 NOR2X1_441 ( .A(_4181_), .B(_4178_), .Y(_4182_) );
	NAND2X1 NAND2X1_762 ( .A(_4174_), .B(_4182_), .Y(_4183_) );
	NOR3X1 NOR3X1_318 ( .A(_4167_), .B(_4152_), .C(_4183_), .Y(_4184_) );
	AOI22X1 AOI22X1_590 ( .A(_3990_), .B(wData[42]), .C(wData[38]), .D(_3992_), .Y(_4185_) );
	AOI22X1 AOI22X1_591 ( .A(_3987_), .B(wData[46]), .C(_3994_), .D(wData[2]), .Y(_4186_) );
	NAND2X1 NAND2X1_763 ( .A(_4185_), .B(_4186_), .Y(_4187_) );
	AOI21X1 AOI21X1_87 ( .A(wData[34]), .B(_3980_), .C(_4187_), .Y(_4188_) );
	INVX1 INVX1_477 ( .A(wData[50]), .Y(_4189_) );
	AOI22X1 AOI22X1_592 ( .A(_4000_), .B(wData[10]), .C(wData[14]), .D(_4001_), .Y(_4190_) );
	OAI21X1 OAI21X1_125 ( .A(_4189_), .B(_3999_), .C(_4190_), .Y(_4191_) );
	AOI22X1 AOI22X1_593 ( .A(_3963_), .B(wData[22]), .C(wData[18]), .D(_3966_), .Y(_4192_) );
	NAND2X1 NAND2X1_764 ( .A(wData[26]), .B(_3970_), .Y(_4193_) );
	AOI22X1 AOI22X1_594 ( .A(_3976_), .B(wData[30]), .C(wData[6]), .D(_3974_), .Y(_4194_) );
	NAND3X1 NAND3X1_183 ( .A(_4193_), .B(_4194_), .C(_4192_), .Y(_4195_) );
	NOR2X1 NOR2X1_442 ( .A(_4191_), .B(_4195_), .Y(_4196_) );
	NAND2X1 NAND2X1_765 ( .A(wData[58]), .B(_3983_), .Y(_4197_) );
	NAND2X1 NAND2X1_766 ( .A(wData[54]), .B(_3984_), .Y(_4198_) );
	NAND2X1 NAND2X1_767 ( .A(_4197_), .B(_4198_), .Y(_4199_) );
	AOI21X1 AOI21X1_88 ( .A(wData[62]), .B(_3986_), .C(_4199_), .Y(_4200_) );
	NAND3X1 NAND3X1_184 ( .A(_4188_), .B(_4200_), .C(_4196_), .Y(_4201_) );
	NOR2X1 NOR2X1_443 ( .A(_3768_), .B(_4201_), .Y(_4202_) );
	AOI21X1 AOI21X1_89 ( .A(_4130_), .B(_4184_), .C(_4202_), .Y(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_2_) );
	AOI21X1 AOI21X1_90 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_4012_), .C(_3769_), .Y(_4203_) );
	AOI22X1 AOI22X1_595 ( .A(_3784_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_4104_), .Y(_4204_) );
	AOI22X1 AOI22X1_596 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_4106_), .C(_3862_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_4205_) );
	NAND3X1 NAND3X1_185 ( .A(_4205_), .B(_4203_), .C(_4204_), .Y(_4206_) );
	AOI22X1 AOI22X1_597 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_3811_), .C(_3809_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_4207_) );
	AOI22X1 AOI22X1_598 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_3882_), .C(_4007_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_4208_) );
	INVX1 INVX1_478 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_4209_) );
	INVX1 INVX1_479 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_4210_) );
	OAI22X1 OAI22X1_102 ( .A(_4209_), .B(_3824_), .C(_3873_), .D(_4210_), .Y(_4211_) );
	INVX1 INVX1_480 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_4212_) );
	NAND2X1 NAND2X1_768 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_3925_), .Y(_4213_) );
	OAI21X1 OAI21X1_126 ( .A(_4212_), .B(_3830_), .C(_4213_), .Y(_4214_) );
	NOR2X1 NOR2X1_444 ( .A(_4211_), .B(_4214_), .Y(_4215_) );
	NAND3X1 NAND3X1_186 ( .A(_4207_), .B(_4208_), .C(_4215_), .Y(_4216_) );
	AND2X2 AND2X2_82 ( .A(_3838_), .B(_3772_), .Y(_4217_) );
	AOI22X1 AOI22X1_599 ( .A(_3777_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_4217_), .Y(_4218_) );
	AND2X2 AND2X2_83 ( .A(_3836_), .B(_3801_), .Y(_4219_) );
	AND2X2 AND2X2_84 ( .A(_3844_), .B(_3801_), .Y(_4220_) );
	AOI22X1 AOI22X1_600 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_4220_), .C(_4219_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_4221_) );
	NAND2X1 NAND2X1_769 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_3929_), .Y(_4222_) );
	NAND2X1 NAND2X1_770 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_3902_), .Y(_4223_) );
	NAND2X1 NAND2X1_771 ( .A(_4222_), .B(_4223_), .Y(_4224_) );
	INVX1 INVX1_481 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_4225_) );
	NAND2X1 NAND2X1_772 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_3901_), .Y(_4226_) );
	OAI21X1 OAI21X1_127 ( .A(_4225_), .B(_3854_), .C(_4226_), .Y(_4227_) );
	NOR2X1 NOR2X1_445 ( .A(_4224_), .B(_4227_), .Y(_4228_) );
	NAND3X1 NAND3X1_187 ( .A(_4218_), .B(_4221_), .C(_4228_), .Y(_4229_) );
	NOR3X1 NOR3X1_319 ( .A(_4216_), .B(_4206_), .C(_4229_), .Y(_4230_) );
	INVX1 INVX1_482 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_4231_) );
	NAND2X1 NAND2X1_773 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_3817_), .Y(_4232_) );
	OAI21X1 OAI21X1_128 ( .A(_3822_), .B(_4231_), .C(_4232_), .Y(_4233_) );
	AOI21X1 AOI21X1_91 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_3797_), .C(_4233_), .Y(_4234_) );
	INVX1 INVX1_483 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_4235_) );
	INVX1 INVX1_484 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_4236_) );
	OAI22X1 OAI22X1_103 ( .A(_4141_), .B(_4236_), .C(_4235_), .D(_3792_), .Y(_4237_) );
	INVX1 INVX1_485 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_4238_) );
	NAND2X1 NAND2X1_774 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_3937_), .Y(_4239_) );
	OAI21X1 OAI21X1_129 ( .A(_3802_), .B(_4238_), .C(_4239_), .Y(_4240_) );
	NOR2X1 NOR2X1_446 ( .A(_4240_), .B(_4237_), .Y(_4241_) );
	INVX1 INVX1_486 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_4242_) );
	INVX1 INVX1_487 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_4243_) );
	OAI22X1 OAI22X1_104 ( .A(_3889_), .B(_4243_), .C(_4242_), .D(_3890_), .Y(_4244_) );
	INVX1 INVX1_488 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_4245_) );
	NAND2X1 NAND2X1_775 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_3936_), .Y(_4246_) );
	OAI21X1 OAI21X1_130 ( .A(_4245_), .B(_3872_), .C(_4246_), .Y(_4247_) );
	NOR2X1 NOR2X1_447 ( .A(_4247_), .B(_4244_), .Y(_4248_) );
	NAND3X1 NAND3X1_188 ( .A(_4234_), .B(_4248_), .C(_4241_), .Y(_4249_) );
	AOI22X1 AOI22X1_601 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_3894_), .C(_3895_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_4250_) );
	AOI22X1 AOI22X1_602 ( .A(_3897_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_3898_), .Y(_4251_) );
	NAND2X1 NAND2X1_776 ( .A(_4250_), .B(_4251_), .Y(_4252_) );
	AOI22X1 AOI22X1_603 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_3905_), .C(_3904_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_4253_) );
	AOI22X1 AOI22X1_604 ( .A(_3848_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_3855_), .Y(_4254_) );
	NAND2X1 NAND2X1_777 ( .A(_4253_), .B(_4254_), .Y(_4255_) );
	NOR2X1 NOR2X1_448 ( .A(_4252_), .B(_4255_), .Y(_4256_) );
	AOI22X1 AOI22X1_605 ( .A(_3909_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_3910_), .Y(_4257_) );
	AOI22X1 AOI22X1_606 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_4145_), .C(_3912_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_4258_) );
	NAND2X1 NAND2X1_778 ( .A(_4258_), .B(_4257_), .Y(_4259_) );
	AOI22X1 AOI22X1_607 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_3916_), .C(_3917_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_4260_) );
	AOI22X1 AOI22X1_608 ( .A(_3919_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_3920_), .Y(_4261_) );
	NAND2X1 NAND2X1_779 ( .A(_4261_), .B(_4260_), .Y(_4262_) );
	NOR2X1 NOR2X1_449 ( .A(_4259_), .B(_4262_), .Y(_4263_) );
	NAND2X1 NAND2X1_780 ( .A(_4263_), .B(_4256_), .Y(_4264_) );
	AOI22X1 AOI22X1_609 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_3926_), .C(_3827_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_4265_) );
	AOI22X1 AOI22X1_610 ( .A(_3850_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_3928_), .Y(_4266_) );
	NAND2X1 NAND2X1_781 ( .A(_4265_), .B(_4266_), .Y(_4267_) );
	AOI22X1 AOI22X1_611 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_3934_), .C(_3932_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_4268_) );
	AOI22X1 AOI22X1_612 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_3864_), .C(_3913_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_4269_) );
	NAND2X1 NAND2X1_782 ( .A(_4269_), .B(_4268_), .Y(_4270_) );
	NOR2X1 NOR2X1_450 ( .A(_4270_), .B(_4267_), .Y(_4271_) );
	AOI22X1 AOI22X1_613 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_3941_), .C(_3942_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_4272_) );
	NAND2X1 NAND2X1_783 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_3944_), .Y(_4273_) );
	NAND2X1 NAND2X1_784 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_3946_), .Y(_4274_) );
	NAND3X1 NAND3X1_189 ( .A(_4273_), .B(_4274_), .C(_4272_), .Y(_4275_) );
	AOI22X1 AOI22X1_614 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_3950_), .C(_3949_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_4276_) );
	AOI22X1 AOI22X1_615 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_3953_), .C(_3952_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_4277_) );
	NAND2X1 NAND2X1_785 ( .A(_4276_), .B(_4277_), .Y(_4278_) );
	NOR2X1 NOR2X1_451 ( .A(_4278_), .B(_4275_), .Y(_4279_) );
	NAND2X1 NAND2X1_786 ( .A(_4271_), .B(_4279_), .Y(_4280_) );
	NOR3X1 NOR3X1_320 ( .A(_4264_), .B(_4249_), .C(_4280_), .Y(_4281_) );
	NAND2X1 NAND2X1_787 ( .A(wData[59]), .B(_3983_), .Y(_4282_) );
	OAI21X1 OAI21X1_131 ( .A(_3767_), .B(wBusy_bF_buf2), .C(_4282_), .Y(_4283_) );
	NAND2X1 NAND2X1_788 ( .A(wData[7]), .B(_3974_), .Y(_4284_) );
	NAND2X1 NAND2X1_789 ( .A(wData[55]), .B(_3984_), .Y(_4285_) );
	AOI22X1 AOI22X1_616 ( .A(wData[63]), .B(_3986_), .C(_3976_), .D(wData[31]), .Y(_4286_) );
	NAND3X1 NAND3X1_190 ( .A(_4284_), .B(_4285_), .C(_4286_), .Y(_4287_) );
	OR2X2 OR2X2_43 ( .A(_4287_), .B(_4283_), .Y(_4288_) );
	INVX1 INVX1_489 ( .A(wData[51]), .Y(_4289_) );
	NAND2X1 NAND2X1_790 ( .A(wData[47]), .B(_3987_), .Y(_4290_) );
	OAI21X1 OAI21X1_132 ( .A(_4289_), .B(_3999_), .C(_4290_), .Y(_4291_) );
	AOI21X1 AOI21X1_92 ( .A(wData[3]), .B(_3994_), .C(_4291_), .Y(_4292_) );
	AOI22X1 AOI22X1_617 ( .A(_4000_), .B(wData[11]), .C(wData[15]), .D(_4001_), .Y(_4293_) );
	AOI22X1 AOI22X1_618 ( .A(_3963_), .B(wData[23]), .C(wData[27]), .D(_3970_), .Y(_4294_) );
	AND2X2 AND2X2_85 ( .A(_4293_), .B(_4294_), .Y(_4295_) );
	NAND2X1 NAND2X1_791 ( .A(wData[39]), .B(_3992_), .Y(_4296_) );
	NAND2X1 NAND2X1_792 ( .A(wData[43]), .B(_3990_), .Y(_4297_) );
	NAND2X1 NAND2X1_793 ( .A(_4296_), .B(_4297_), .Y(_4298_) );
	NAND2X1 NAND2X1_794 ( .A(wData[19]), .B(_3966_), .Y(_4299_) );
	NAND2X1 NAND2X1_795 ( .A(wData[35]), .B(_3980_), .Y(_4300_) );
	NAND2X1 NAND2X1_796 ( .A(_4299_), .B(_4300_), .Y(_4301_) );
	NOR2X1 NOR2X1_452 ( .A(_4298_), .B(_4301_), .Y(_4302_) );
	NAND3X1 NAND3X1_191 ( .A(_4295_), .B(_4292_), .C(_4302_), .Y(_4303_) );
	NOR2X1 NOR2X1_453 ( .A(_4288_), .B(_4303_), .Y(_4304_) );
	AOI21X1 AOI21X1_93 ( .A(_4230_), .B(_4281_), .C(_4304_), .Y(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_3_) );
	INVX1 INVX1_490 ( .A(wSelec[88]), .Y(_4305_) );
	NOR2X1 NOR2X1_454 ( .A(wBusy_bF_buf1), .B(_4305_), .Y(_4306_) );
	INVX1 INVX1_491 ( .A(_4306_), .Y(_4307_) );
	INVX1 INVX1_492 ( .A(wSelec[98]), .Y(_4308_) );
	NAND2X1 NAND2X1_797 ( .A(wSelec[97]), .B(_4308_), .Y(_4309_) );
	INVX2 INVX2_13 ( .A(_4309_), .Y(_4310_) );
	OR2X2 OR2X2_44 ( .A(wSelec[94]), .B(wSelec[93]), .Y(_4311_) );
	INVX1 INVX1_493 ( .A(wSelec[96]), .Y(_4312_) );
	NAND2X1 NAND2X1_798 ( .A(wSelec[95]), .B(_4312_), .Y(_4313_) );
	NOR2X1 NOR2X1_455 ( .A(_4311_), .B(_4313_), .Y(_4314_) );
	AND2X2 AND2X2_86 ( .A(_4314_), .B(_4310_), .Y(_4315_) );
	AOI21X1 AOI21X1_94 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_4315_), .C(_4307_), .Y(_4316_) );
	INVX1 INVX1_494 ( .A(wSelec[94]), .Y(_4317_) );
	NAND2X1 NAND2X1_799 ( .A(wSelec[93]), .B(_4317_), .Y(_4318_) );
	OR2X2 OR2X2_45 ( .A(wSelec[95]), .B(wSelec[96]), .Y(_4319_) );
	NOR2X1 NOR2X1_456 ( .A(_4319_), .B(_4318_), .Y(_4320_) );
	NAND2X1 NAND2X1_800 ( .A(_4310_), .B(_4320_), .Y(_4321_) );
	INVX1 INVX1_495 ( .A(_4321_), .Y(_4322_) );
	INVX1 INVX1_496 ( .A(wSelec[93]), .Y(_4323_) );
	NAND2X1 NAND2X1_801 ( .A(wSelec[94]), .B(_4323_), .Y(_4324_) );
	INVX1 INVX1_497 ( .A(wSelec[95]), .Y(_4325_) );
	NAND2X1 NAND2X1_802 ( .A(wSelec[96]), .B(_4325_), .Y(_4326_) );
	NOR2X1 NOR2X1_457 ( .A(_4324_), .B(_4326_), .Y(_4327_) );
	NAND2X1 NAND2X1_803 ( .A(wSelec[97]), .B(wSelec[98]), .Y(_4328_) );
	INVX1 INVX1_498 ( .A(_4328_), .Y(_4329_) );
	NAND2X1 NAND2X1_804 ( .A(_4329_), .B(_4327_), .Y(_4330_) );
	INVX1 INVX1_499 ( .A(_4330_), .Y(_4331_) );
	AOI22X1 AOI22X1_619 ( .A(_4322_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_4331_), .Y(_4332_) );
	OR2X2 OR2X2_46 ( .A(_4318_), .B(_4319_), .Y(_4333_) );
	OR2X2 OR2X2_47 ( .A(wSelec[97]), .B(wSelec[98]), .Y(_4334_) );
	NOR2X1 NOR2X1_458 ( .A(_4334_), .B(_4333_), .Y(_4335_) );
	NOR2X1 NOR2X1_459 ( .A(_4313_), .B(_4318_), .Y(_4336_) );
	INVX1 INVX1_500 ( .A(wSelec[97]), .Y(_4337_) );
	NAND2X1 NAND2X1_805 ( .A(wSelec[98]), .B(_4337_), .Y(_4338_) );
	INVX2 INVX2_14 ( .A(_4338_), .Y(_4339_) );
	NAND2X1 NAND2X1_806 ( .A(_4339_), .B(_4336_), .Y(_4340_) );
	INVX1 INVX1_501 ( .A(_4340_), .Y(_4341_) );
	AOI22X1 AOI22X1_620 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_4335_), .C(_4341_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_4342_) );
	NAND3X1 NAND3X1_192 ( .A(_4316_), .B(_4342_), .C(_4332_), .Y(_4343_) );
	NOR2X1 NOR2X1_460 ( .A(wSelec[94]), .B(wSelec[93]), .Y(_4344_) );
	NOR2X1 NOR2X1_461 ( .A(wSelec[95]), .B(wSelec[96]), .Y(_4345_) );
	NAND2X1 NAND2X1_807 ( .A(_4344_), .B(_4345_), .Y(_4346_) );
	NOR2X1 NOR2X1_462 ( .A(_4309_), .B(_4346_), .Y(_4347_) );
	NAND2X1 NAND2X1_808 ( .A(wSelec[94]), .B(wSelec[93]), .Y(_4348_) );
	NOR3X1 NOR3X1_321 ( .A(_4319_), .B(_4348_), .C(_4309_), .Y(_4349_) );
	AOI22X1 AOI22X1_621 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_4349_), .C(_4347_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_4350_) );
	INVX1 INVX1_502 ( .A(_4334_), .Y(_4351_) );
	NOR2X1 NOR2X1_463 ( .A(_4319_), .B(_4324_), .Y(_4352_) );
	AND2X2 AND2X2_87 ( .A(_4352_), .B(_4351_), .Y(_4353_) );
	NAND2X1 NAND2X1_809 ( .A(wSelec[95]), .B(wSelec[96]), .Y(_4354_) );
	NOR3X1 NOR3X1_322 ( .A(_4328_), .B(_4348_), .C(_4354_), .Y(_4355_) );
	AOI22X1 AOI22X1_622 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_4355_), .C(_4353_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_4356_) );
	INVX1 INVX1_503 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_4357_) );
	INVX1 INVX1_504 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_4358_) );
	NOR2X1 NOR2X1_464 ( .A(_4318_), .B(_4326_), .Y(_4359_) );
	NAND2X1 NAND2X1_810 ( .A(_4329_), .B(_4359_), .Y(_4360_) );
	NOR2X1 NOR2X1_465 ( .A(_4348_), .B(_4354_), .Y(_4361_) );
	NAND2X1 NAND2X1_811 ( .A(_4361_), .B(_4339_), .Y(_4362_) );
	OAI22X1 OAI22X1_105 ( .A(_4357_), .B(_4362_), .C(_4360_), .D(_4358_), .Y(_4363_) );
	INVX1 INVX1_505 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_4364_) );
	NOR3X1 NOR3X1_323 ( .A(_4309_), .B(_4324_), .C(_4326_), .Y(_4365_) );
	NAND2X1 NAND2X1_812 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_4365_), .Y(_4366_) );
	NOR2X1 NOR2X1_466 ( .A(_4348_), .B(_4313_), .Y(_4367_) );
	NAND2X1 NAND2X1_813 ( .A(_4339_), .B(_4367_), .Y(_4368_) );
	OAI21X1 OAI21X1_133 ( .A(_4364_), .B(_4368_), .C(_4366_), .Y(_4369_) );
	NOR2X1 NOR2X1_467 ( .A(_4363_), .B(_4369_), .Y(_4370_) );
	NAND3X1 NAND3X1_193 ( .A(_4350_), .B(_4356_), .C(_4370_), .Y(_4371_) );
	INVX1 INVX1_506 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_4372_) );
	INVX1 INVX1_507 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_4373_) );
	NOR2X1 NOR2X1_468 ( .A(_4313_), .B(_4324_), .Y(_4374_) );
	NAND2X1 NAND2X1_814 ( .A(_4310_), .B(_4374_), .Y(_4375_) );
	NOR2X1 NOR2X1_469 ( .A(_4311_), .B(_4326_), .Y(_4376_) );
	NAND2X1 NAND2X1_815 ( .A(_4310_), .B(_4376_), .Y(_4377_) );
	OAI22X1 OAI22X1_106 ( .A(_4377_), .B(_4372_), .C(_4373_), .D(_4375_), .Y(_4378_) );
	INVX1 INVX1_508 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_4379_) );
	INVX1 INVX1_509 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_4380_) );
	NAND2X1 NAND2X1_816 ( .A(_4339_), .B(_4374_), .Y(_4381_) );
	NOR2X1 NOR2X1_470 ( .A(_4348_), .B(_4319_), .Y(_4382_) );
	NAND2X1 NAND2X1_817 ( .A(_4339_), .B(_4382_), .Y(_4383_) );
	OAI22X1 OAI22X1_107 ( .A(_4379_), .B(_4383_), .C(_4381_), .D(_4380_), .Y(_4384_) );
	NOR2X1 NOR2X1_471 ( .A(_4384_), .B(_4378_), .Y(_4385_) );
	NOR3X1 NOR3X1_324 ( .A(_4318_), .B(_4354_), .C(_4338_), .Y(_4386_) );
	NAND2X1 NAND2X1_818 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_4386_), .Y(_4387_) );
	NOR3X1 NOR3X1_325 ( .A(_4326_), .B(_4348_), .C(_4338_), .Y(_4388_) );
	NAND2X1 NAND2X1_819 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_4388_), .Y(_4389_) );
	NAND2X1 NAND2X1_820 ( .A(_4387_), .B(_4389_), .Y(_4390_) );
	INVX1 INVX1_510 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_4391_) );
	NAND2X1 NAND2X1_821 ( .A(_4329_), .B(_4314_), .Y(_4392_) );
	NOR3X1 NOR3X1_326 ( .A(_4324_), .B(_4326_), .C(_4338_), .Y(_4393_) );
	NAND2X1 NAND2X1_822 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_4393_), .Y(_4394_) );
	OAI21X1 OAI21X1_134 ( .A(_4391_), .B(_4392_), .C(_4394_), .Y(_4395_) );
	NOR2X1 NOR2X1_472 ( .A(_4390_), .B(_4395_), .Y(_4396_) );
	NAND2X1 NAND2X1_823 ( .A(_4385_), .B(_4396_), .Y(_4397_) );
	NOR3X1 NOR3X1_327 ( .A(_4343_), .B(_4397_), .C(_4371_), .Y(_4398_) );
	NAND2X1 NAND2X1_824 ( .A(_4310_), .B(_4367_), .Y(_4399_) );
	INVX1 INVX1_511 ( .A(_4399_), .Y(_4400_) );
	INVX1 INVX1_512 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_4401_) );
	NOR3X1 NOR3X1_328 ( .A(_4311_), .B(_4334_), .C(_4313_), .Y(_4402_) );
	NAND2X1 NAND2X1_825 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_4402_), .Y(_4403_) );
	NAND2X1 NAND2X1_826 ( .A(_4351_), .B(_4374_), .Y(_4404_) );
	OAI21X1 OAI21X1_135 ( .A(_4404_), .B(_4401_), .C(_4403_), .Y(_4405_) );
	AOI21X1 AOI21X1_95 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_4400_), .C(_4405_), .Y(_4406_) );
	INVX1 INVX1_513 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_4407_) );
	INVX1 INVX1_514 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_4408_) );
	NOR2X1 NOR2X1_473 ( .A(_4354_), .B(_4311_), .Y(_4409_) );
	NAND2X1 NAND2X1_827 ( .A(_4310_), .B(_4409_), .Y(_4410_) );
	NAND2X1 NAND2X1_828 ( .A(_4351_), .B(_4336_), .Y(_4411_) );
	OAI22X1 OAI22X1_108 ( .A(_4408_), .B(_4410_), .C(_4411_), .D(_4407_), .Y(_4412_) );
	INVX1 INVX1_515 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_4413_) );
	INVX1 INVX1_516 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_4414_) );
	NAND2X1 NAND2X1_829 ( .A(_4310_), .B(_4336_), .Y(_4415_) );
	NAND2X1 NAND2X1_830 ( .A(_4351_), .B(_4382_), .Y(_4416_) );
	OAI22X1 OAI22X1_109 ( .A(_4413_), .B(_4416_), .C(_4415_), .D(_4414_), .Y(_4417_) );
	NOR2X1 NOR2X1_474 ( .A(_4412_), .B(_4417_), .Y(_4418_) );
	INVX1 INVX1_517 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_4419_) );
	NOR3X1 NOR3X1_329 ( .A(_4334_), .B(_4348_), .C(_4313_), .Y(_4420_) );
	NAND2X1 NAND2X1_831 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_4420_), .Y(_4421_) );
	OR2X2 OR2X2_48 ( .A(_4346_), .B(_4328_), .Y(_4422_) );
	OAI21X1 OAI21X1_136 ( .A(_4419_), .B(_4422_), .C(_4421_), .Y(_4423_) );
	INVX1 INVX1_518 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_4424_) );
	INVX1 INVX1_519 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_4425_) );
	NOR2X1 NOR2X1_475 ( .A(_4354_), .B(_4324_), .Y(_4426_) );
	NAND2X1 NAND2X1_832 ( .A(_4310_), .B(_4426_), .Y(_4427_) );
	NAND2X1 NAND2X1_833 ( .A(_4329_), .B(_4320_), .Y(_4428_) );
	OAI22X1 OAI22X1_110 ( .A(_4427_), .B(_4425_), .C(_4424_), .D(_4428_), .Y(_4429_) );
	NOR2X1 NOR2X1_476 ( .A(_4423_), .B(_4429_), .Y(_4430_) );
	NAND3X1 NAND3X1_194 ( .A(_4406_), .B(_4430_), .C(_4418_), .Y(_4431_) );
	NOR3X1 NOR3X1_330 ( .A(_4311_), .B(_4319_), .C(_4334_), .Y(_4432_) );
	NOR3X1 NOR3X1_331 ( .A(_4328_), .B(_4354_), .C(_4318_), .Y(_4433_) );
	AOI22X1 AOI22X1_623 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_4432_), .C(_4433_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_4434_) );
	NOR3X1 NOR3X1_332 ( .A(_4328_), .B(_4354_), .C(_4324_), .Y(_4435_) );
	NOR3X1 NOR3X1_333 ( .A(_4328_), .B(_4348_), .C(_4326_), .Y(_4436_) );
	AOI22X1 AOI22X1_624 ( .A(_4435_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_4436_), .Y(_4437_) );
	NAND2X1 NAND2X1_834 ( .A(_4434_), .B(_4437_), .Y(_4438_) );
	NOR3X1 NOR3X1_334 ( .A(_4326_), .B(_4311_), .C(_4338_), .Y(_4439_) );
	NOR3X1 NOR3X1_335 ( .A(_4318_), .B(_4326_), .C(_4338_), .Y(_4440_) );
	AOI22X1 AOI22X1_625 ( .A(_4439_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_4440_), .Y(_4441_) );
	NOR3X1 NOR3X1_336 ( .A(_4309_), .B(_4354_), .C(_4318_), .Y(_4442_) );
	NOR3X1 NOR3X1_337 ( .A(_4348_), .B(_4354_), .C(_4309_), .Y(_4443_) );
	AOI22X1 AOI22X1_626 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_4443_), .C(_4442_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_4444_) );
	NAND2X1 NAND2X1_835 ( .A(_4444_), .B(_4441_), .Y(_4445_) );
	NOR2X1 NOR2X1_477 ( .A(_4438_), .B(_4445_), .Y(_4446_) );
	NOR3X1 NOR3X1_338 ( .A(_4334_), .B(_4354_), .C(_4318_), .Y(_4447_) );
	NOR3X1 NOR3X1_339 ( .A(_4334_), .B(_4354_), .C(_4324_), .Y(_4448_) );
	AOI22X1 AOI22X1_627 ( .A(_4447_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_4448_), .Y(_4449_) );
	NOR3X1 NOR3X1_340 ( .A(_4334_), .B(_4348_), .C(_4326_), .Y(_4450_) );
	NOR3X1 NOR3X1_341 ( .A(_4309_), .B(_4319_), .C(_4324_), .Y(_4451_) );
	AOI22X1 AOI22X1_628 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_4450_), .C(_4451_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_4452_) );
	NAND2X1 NAND2X1_836 ( .A(_4449_), .B(_4452_), .Y(_4453_) );
	NOR3X1 NOR3X1_342 ( .A(_4348_), .B(_4354_), .C(_4334_), .Y(_4454_) );
	NOR3X1 NOR3X1_343 ( .A(_4324_), .B(_4319_), .C(_4338_), .Y(_4455_) );
	AOI22X1 AOI22X1_629 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_4454_), .C(_4455_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_4456_) );
	NOR3X1 NOR3X1_344 ( .A(_4311_), .B(_4319_), .C(_4338_), .Y(_4457_) );
	NOR3X1 NOR3X1_345 ( .A(_4311_), .B(_4354_), .C(_4338_), .Y(_4458_) );
	AOI22X1 AOI22X1_630 ( .A(_4457_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_4458_), .Y(_4459_) );
	NAND2X1 NAND2X1_837 ( .A(_4459_), .B(_4456_), .Y(_4460_) );
	NOR2X1 NOR2X1_478 ( .A(_4453_), .B(_4460_), .Y(_4461_) );
	NAND2X1 NAND2X1_838 ( .A(_4461_), .B(_4446_), .Y(_4462_) );
	NOR3X1 NOR3X1_346 ( .A(_4309_), .B(_4348_), .C(_4326_), .Y(_4463_) );
	NOR3X1 NOR3X1_347 ( .A(_4319_), .B(_4328_), .C(_4324_), .Y(_4464_) );
	AOI22X1 AOI22X1_631 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_4464_), .C(_4463_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_4465_) );
	NOR3X1 NOR3X1_348 ( .A(_4313_), .B(_4311_), .C(_4338_), .Y(_4466_) );
	NOR3X1 NOR3X1_349 ( .A(_4324_), .B(_4354_), .C(_4338_), .Y(_4467_) );
	AOI22X1 AOI22X1_632 ( .A(_4466_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_4467_), .Y(_4468_) );
	NAND2X1 NAND2X1_839 ( .A(_4465_), .B(_4468_), .Y(_4469_) );
	NOR3X1 NOR3X1_350 ( .A(_4309_), .B(_4318_), .C(_4326_), .Y(_4470_) );
	NAND2X1 NAND2X1_840 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_4470_), .Y(_4471_) );
	NOR3X1 NOR3X1_351 ( .A(_4328_), .B(_4348_), .C(_4313_), .Y(_4472_) );
	NAND2X1 NAND2X1_841 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_4472_), .Y(_4473_) );
	NOR3X1 NOR3X1_352 ( .A(_4311_), .B(_4354_), .C(_4334_), .Y(_4474_) );
	NOR3X1 NOR3X1_353 ( .A(_4311_), .B(_4328_), .C(_4326_), .Y(_4475_) );
	AOI22X1 AOI22X1_633 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_4474_), .C(_4475_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_4476_) );
	NAND3X1 NAND3X1_195 ( .A(_4471_), .B(_4473_), .C(_4476_), .Y(_4477_) );
	NOR2X1 NOR2X1_479 ( .A(_4477_), .B(_4469_), .Y(_4478_) );
	NOR3X1 NOR3X1_354 ( .A(_4311_), .B(_4334_), .C(_4326_), .Y(_4479_) );
	NOR3X1 NOR3X1_355 ( .A(_4313_), .B(_4328_), .C(_4318_), .Y(_4480_) );
	AOI22X1 AOI22X1_634 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_4479_), .C(_4480_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_4481_) );
	NOR3X1 NOR3X1_356 ( .A(_4313_), .B(_4328_), .C(_4324_), .Y(_4482_) );
	NAND2X1 NAND2X1_842 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_4482_), .Y(_4483_) );
	NOR3X1 NOR3X1_357 ( .A(_4318_), .B(_4319_), .C(_4338_), .Y(_4484_) );
	NAND2X1 NAND2X1_843 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_4484_), .Y(_4485_) );
	NAND3X1 NAND3X1_196 ( .A(_4483_), .B(_4485_), .C(_4481_), .Y(_4486_) );
	NOR3X1 NOR3X1_358 ( .A(_4318_), .B(_4334_), .C(_4326_), .Y(_4487_) );
	NOR3X1 NOR3X1_359 ( .A(_4328_), .B(_4354_), .C(_4311_), .Y(_4488_) );
	AOI22X1 AOI22X1_635 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_4488_), .C(_4487_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_4489_) );
	NOR3X1 NOR3X1_360 ( .A(_4324_), .B(_4334_), .C(_4326_), .Y(_4490_) );
	NOR3X1 NOR3X1_361 ( .A(_4328_), .B(_4348_), .C(_4319_), .Y(_4491_) );
	AOI22X1 AOI22X1_636 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_4491_), .C(_4490_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_4492_) );
	NAND2X1 NAND2X1_844 ( .A(_4489_), .B(_4492_), .Y(_4493_) );
	NOR2X1 NOR2X1_480 ( .A(_4493_), .B(_4486_), .Y(_4494_) );
	NAND2X1 NAND2X1_845 ( .A(_4478_), .B(_4494_), .Y(_4495_) );
	NOR3X1 NOR3X1_362 ( .A(_4462_), .B(_4431_), .C(_4495_), .Y(_4496_) );
	INVX1 INVX1_520 ( .A(wSelec[90]), .Y(_4497_) );
	NAND2X1 NAND2X1_846 ( .A(wSelec[89]), .B(_4497_), .Y(_4498_) );
	INVX1 INVX1_521 ( .A(wSelec[92]), .Y(_4499_) );
	NAND2X1 NAND2X1_847 ( .A(wSelec[91]), .B(_4499_), .Y(_4500_) );
	NOR2X1 NOR2X1_481 ( .A(_4498_), .B(_4500_), .Y(_4501_) );
	NOR2X1 NOR2X1_482 ( .A(wSelec[90]), .B(wSelec[89]), .Y(_4502_) );
	INVX1 INVX1_522 ( .A(_4502_), .Y(_4503_) );
	NOR2X1 NOR2X1_483 ( .A(_4500_), .B(_4503_), .Y(_4504_) );
	AOI22X1 AOI22X1_637 ( .A(wData[20]), .B(_4501_), .C(_4504_), .D(wData[16]), .Y(_4505_) );
	INVX1 INVX1_523 ( .A(wSelec[89]), .Y(_4506_) );
	NAND2X1 NAND2X1_848 ( .A(wSelec[90]), .B(_4506_), .Y(_4507_) );
	NOR2X1 NOR2X1_484 ( .A(_4507_), .B(_4500_), .Y(_4508_) );
	NAND2X1 NAND2X1_849 ( .A(wData[24]), .B(_4508_), .Y(_4509_) );
	INVX1 INVX1_524 ( .A(wSelec[91]), .Y(_4510_) );
	NAND2X1 NAND2X1_850 ( .A(_4510_), .B(_4499_), .Y(_4511_) );
	NOR2X1 NOR2X1_485 ( .A(_4498_), .B(_4511_), .Y(_4512_) );
	NAND2X1 NAND2X1_851 ( .A(wSelec[90]), .B(wSelec[89]), .Y(_4513_) );
	NOR2X1 NOR2X1_486 ( .A(_4513_), .B(_4500_), .Y(_4514_) );
	AOI22X1 AOI22X1_638 ( .A(_4514_), .B(wData[28]), .C(wData[4]), .D(_4512_), .Y(_4515_) );
	NAND3X1 NAND3X1_197 ( .A(_4509_), .B(_4515_), .C(_4505_), .Y(_4516_) );
	NAND2X1 NAND2X1_852 ( .A(wSelec[92]), .B(_4510_), .Y(_4517_) );
	NOR2X1 NOR2X1_487 ( .A(_4517_), .B(_4503_), .Y(_4518_) );
	NAND2X1 NAND2X1_853 ( .A(wData[32]), .B(_4518_), .Y(_4519_) );
	NAND2X1 NAND2X1_854 ( .A(wSelec[91]), .B(wSelec[92]), .Y(_4520_) );
	NOR2X1 NOR2X1_488 ( .A(_4520_), .B(_4507_), .Y(_4521_) );
	NOR2X1 NOR2X1_489 ( .A(_4520_), .B(_4498_), .Y(_4522_) );
	AOI22X1 AOI22X1_639 ( .A(_4521_), .B(wData[56]), .C(wData[52]), .D(_4522_), .Y(_4523_) );
	NOR2X1 NOR2X1_490 ( .A(_4513_), .B(_4520_), .Y(_4524_) );
	NOR2X1 NOR2X1_491 ( .A(_4513_), .B(_4517_), .Y(_4525_) );
	AOI22X1 AOI22X1_640 ( .A(wData[60]), .B(_4524_), .C(_4525_), .D(wData[44]), .Y(_4526_) );
	NAND3X1 NAND3X1_198 ( .A(_4519_), .B(_4526_), .C(_4523_), .Y(_4527_) );
	NOR2X1 NOR2X1_492 ( .A(_4507_), .B(_4517_), .Y(_4528_) );
	NAND2X1 NAND2X1_855 ( .A(wData[40]), .B(_4528_), .Y(_4529_) );
	NOR2X1 NOR2X1_493 ( .A(_4517_), .B(_4498_), .Y(_4530_) );
	NAND2X1 NAND2X1_856 ( .A(wData[36]), .B(_4530_), .Y(_4531_) );
	NOR2X1 NOR2X1_494 ( .A(_4511_), .B(_4503_), .Y(_4532_) );
	NAND2X1 NAND2X1_857 ( .A(wData[0]), .B(_4532_), .Y(_4533_) );
	NAND3X1 NAND3X1_199 ( .A(_4529_), .B(_4531_), .C(_4533_), .Y(_4534_) );
	INVX1 INVX1_525 ( .A(wData[48]), .Y(_4535_) );
	NOR2X1 NOR2X1_495 ( .A(_4510_), .B(_4499_), .Y(_4536_) );
	NAND2X1 NAND2X1_858 ( .A(_4502_), .B(_4536_), .Y(_4537_) );
	NOR2X1 NOR2X1_496 ( .A(_4507_), .B(_4511_), .Y(_4538_) );
	NOR2X1 NOR2X1_497 ( .A(_4513_), .B(_4511_), .Y(_4539_) );
	AOI22X1 AOI22X1_641 ( .A(_4538_), .B(wData[8]), .C(wData[12]), .D(_4539_), .Y(_4540_) );
	OAI21X1 OAI21X1_137 ( .A(_4535_), .B(_4537_), .C(_4540_), .Y(_4541_) );
	OR2X2 OR2X2_49 ( .A(_4541_), .B(_4534_), .Y(_4542_) );
	NOR3X1 NOR3X1_363 ( .A(_4516_), .B(_4527_), .C(_4542_), .Y(_4543_) );
	AND2X2 AND2X2_88 ( .A(_4543_), .B(_4307_), .Y(_4544_) );
	AOI21X1 AOI21X1_96 ( .A(_4398_), .B(_4496_), .C(_4544_), .Y(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_0_) );
	INVX1 INVX1_526 ( .A(_4415_), .Y(_4545_) );
	AOI21X1 AOI21X1_97 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_4545_), .C(_4307_), .Y(_4546_) );
	AOI22X1 AOI22X1_642 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_4315_), .C(_4331_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_4547_) );
	AOI22X1 AOI22X1_643 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_4335_), .C(_4341_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_4548_) );
	NAND3X1 NAND3X1_200 ( .A(_4546_), .B(_4547_), .C(_4548_), .Y(_4549_) );
	INVX1 INVX1_527 ( .A(_4375_), .Y(_4550_) );
	AOI22X1 AOI22X1_644 ( .A(_4400_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_4550_), .Y(_4551_) );
	AOI22X1 AOI22X1_645 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_4474_), .C(_4353_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_4552_) );
	INVX1 INVX1_528 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_4553_) );
	INVX1 INVX1_529 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_4554_) );
	OAI22X1 OAI22X1_111 ( .A(_4553_), .B(_4362_), .C(_4360_), .D(_4554_), .Y(_4555_) );
	INVX1 INVX1_530 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_4556_) );
	NAND2X1 NAND2X1_859 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_4463_), .Y(_4557_) );
	OAI21X1 OAI21X1_138 ( .A(_4556_), .B(_4368_), .C(_4557_), .Y(_4558_) );
	NOR2X1 NOR2X1_498 ( .A(_4555_), .B(_4558_), .Y(_4559_) );
	NAND3X1 NAND3X1_201 ( .A(_4551_), .B(_4552_), .C(_4559_), .Y(_4560_) );
	INVX1 INVX1_531 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_4561_) );
	NAND2X1 NAND2X1_860 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_4347_), .Y(_4562_) );
	OAI21X1 OAI21X1_139 ( .A(_4561_), .B(_4377_), .C(_4562_), .Y(_4563_) );
	INVX1 INVX1_532 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_4564_) );
	INVX1 INVX1_533 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_4565_) );
	OAI22X1 OAI22X1_112 ( .A(_4564_), .B(_4383_), .C(_4381_), .D(_4565_), .Y(_4566_) );
	NOR2X1 NOR2X1_499 ( .A(_4566_), .B(_4563_), .Y(_4567_) );
	AOI22X1 AOI22X1_646 ( .A(_4467_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_4440_), .Y(_4568_) );
	AND2X2 AND2X2_89 ( .A(_4314_), .B(_4329_), .Y(_4569_) );
	AOI22X1 AOI22X1_647 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_4439_), .C(_4569_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_4570_) );
	NAND3X1 NAND3X1_202 ( .A(_4568_), .B(_4570_), .C(_4567_), .Y(_4571_) );
	NOR3X1 NOR3X1_364 ( .A(_4571_), .B(_4549_), .C(_4560_), .Y(_4572_) );
	INVX1 INVX1_534 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_4573_) );
	NAND2X1 NAND2X1_861 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_4402_), .Y(_4574_) );
	OAI21X1 OAI21X1_140 ( .A(_4404_), .B(_4573_), .C(_4574_), .Y(_4575_) );
	AOI21X1 AOI21X1_98 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_4451_), .C(_4575_), .Y(_4576_) );
	INVX1 INVX1_535 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_4577_) );
	INVX1 INVX1_536 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_4578_) );
	OAI22X1 OAI22X1_113 ( .A(_4578_), .B(_4410_), .C(_4411_), .D(_4577_), .Y(_4579_) );
	INVX1 INVX1_537 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_4580_) );
	NAND2X1 NAND2X1_862 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_4420_), .Y(_4581_) );
	OAI21X1 OAI21X1_141 ( .A(_4321_), .B(_4580_), .C(_4581_), .Y(_4582_) );
	NOR2X1 NOR2X1_500 ( .A(_4582_), .B(_4579_), .Y(_4583_) );
	INVX1 INVX1_538 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_4584_) );
	INVX1 INVX1_539 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_4585_) );
	OAI22X1 OAI22X1_114 ( .A(_4416_), .B(_4585_), .C(_4422_), .D(_4584_), .Y(_4586_) );
	INVX1 INVX1_540 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_4587_) );
	NOR2X1 NOR2X1_501 ( .A(_4587_), .B(_4427_), .Y(_4588_) );
	INVX1 INVX1_541 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_4589_) );
	NOR2X1 NOR2X1_502 ( .A(_4589_), .B(_4428_), .Y(_4590_) );
	NOR3X1 NOR3X1_365 ( .A(_4588_), .B(_4586_), .C(_4590_), .Y(_4591_) );
	NAND3X1 NAND3X1_203 ( .A(_4583_), .B(_4576_), .C(_4591_), .Y(_4592_) );
	AOI22X1 AOI22X1_648 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_4432_), .C(_4433_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_4593_) );
	AOI22X1 AOI22X1_649 ( .A(_4435_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_4436_), .Y(_4594_) );
	NAND2X1 NAND2X1_863 ( .A(_4593_), .B(_4594_), .Y(_4595_) );
	AOI22X1 AOI22X1_650 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_4443_), .C(_4442_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_4596_) );
	AOI22X1 AOI22X1_651 ( .A(_4386_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_4393_), .Y(_4597_) );
	NAND2X1 NAND2X1_864 ( .A(_4596_), .B(_4597_), .Y(_4598_) );
	NOR2X1 NOR2X1_503 ( .A(_4595_), .B(_4598_), .Y(_4599_) );
	AOI22X1 AOI22X1_652 ( .A(_4447_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_4448_), .Y(_4600_) );
	AOI22X1 AOI22X1_653 ( .A(_4349_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_4450_), .Y(_4601_) );
	NAND2X1 NAND2X1_865 ( .A(_4600_), .B(_4601_), .Y(_4602_) );
	AOI22X1 AOI22X1_654 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_4454_), .C(_4455_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_4603_) );
	AOI22X1 AOI22X1_655 ( .A(_4457_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_4458_), .Y(_4604_) );
	NAND2X1 NAND2X1_866 ( .A(_4604_), .B(_4603_), .Y(_4605_) );
	NOR2X1 NOR2X1_504 ( .A(_4602_), .B(_4605_), .Y(_4606_) );
	NAND2X1 NAND2X1_867 ( .A(_4606_), .B(_4599_), .Y(_4607_) );
	AOI22X1 AOI22X1_656 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_4464_), .C(_4365_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_4608_) );
	AOI22X1 AOI22X1_657 ( .A(_4388_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_4466_), .Y(_4609_) );
	NAND2X1 NAND2X1_868 ( .A(_4608_), .B(_4609_), .Y(_4610_) );
	AOI22X1 AOI22X1_658 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_4355_), .C(_4475_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_4611_) );
	NAND2X1 NAND2X1_869 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_4470_), .Y(_4612_) );
	NAND2X1 NAND2X1_870 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_4472_), .Y(_4613_) );
	NAND3X1 NAND3X1_204 ( .A(_4612_), .B(_4613_), .C(_4611_), .Y(_4614_) );
	NOR2X1 NOR2X1_505 ( .A(_4614_), .B(_4610_), .Y(_4615_) );
	AOI22X1 AOI22X1_659 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_4479_), .C(_4480_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_4616_) );
	NAND2X1 NAND2X1_871 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_4482_), .Y(_4617_) );
	NAND2X1 NAND2X1_872 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_4484_), .Y(_4618_) );
	NAND3X1 NAND3X1_205 ( .A(_4617_), .B(_4618_), .C(_4616_), .Y(_4619_) );
	AOI22X1 AOI22X1_660 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_4488_), .C(_4487_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_4620_) );
	AOI22X1 AOI22X1_661 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_4491_), .C(_4490_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_4621_) );
	NAND2X1 NAND2X1_873 ( .A(_4620_), .B(_4621_), .Y(_4622_) );
	NOR2X1 NOR2X1_506 ( .A(_4622_), .B(_4619_), .Y(_4623_) );
	NAND2X1 NAND2X1_874 ( .A(_4615_), .B(_4623_), .Y(_4624_) );
	NOR3X1 NOR3X1_366 ( .A(_4607_), .B(_4592_), .C(_4624_), .Y(_4625_) );
	AOI21X1 AOI21X1_99 ( .A(wData[21]), .B(_4501_), .C(_4306_), .Y(_4626_) );
	AOI22X1 AOI22X1_662 ( .A(_4504_), .B(wData[17]), .C(wData[1]), .D(_4532_), .Y(_4627_) );
	AOI22X1 AOI22X1_663 ( .A(_4525_), .B(wData[45]), .C(wData[25]), .D(_4508_), .Y(_4628_) );
	NAND3X1 NAND3X1_206 ( .A(_4626_), .B(_4628_), .C(_4627_), .Y(_4629_) );
	NAND3X1 NAND3X1_207 ( .A(wData[49]), .B(_4502_), .C(_4536_), .Y(_4630_) );
	AOI22X1 AOI22X1_664 ( .A(wData[61]), .B(_4524_), .C(_4512_), .D(wData[5]), .Y(_4631_) );
	AND2X2 AND2X2_90 ( .A(_4631_), .B(_4630_), .Y(_4632_) );
	AOI22X1 AOI22X1_665 ( .A(_4521_), .B(wData[57]), .C(wData[41]), .D(_4528_), .Y(_4633_) );
	AOI22X1 AOI22X1_666 ( .A(wData[53]), .B(_4522_), .C(_4518_), .D(wData[33]), .Y(_4634_) );
	AND2X2 AND2X2_91 ( .A(_4634_), .B(_4633_), .Y(_4635_) );
	AOI22X1 AOI22X1_667 ( .A(_4538_), .B(wData[9]), .C(wData[13]), .D(_4539_), .Y(_4636_) );
	AOI22X1 AOI22X1_668 ( .A(_4514_), .B(wData[29]), .C(wData[37]), .D(_4530_), .Y(_4637_) );
	AND2X2 AND2X2_92 ( .A(_4636_), .B(_4637_), .Y(_4638_) );
	NAND3X1 NAND3X1_208 ( .A(_4632_), .B(_4638_), .C(_4635_), .Y(_4639_) );
	NOR2X1 NOR2X1_507 ( .A(_4629_), .B(_4639_), .Y(_4640_) );
	AOI21X1 AOI21X1_100 ( .A(_4572_), .B(_4625_), .C(_4640_), .Y(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_1_) );
	AOI21X1 AOI21X1_101 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_4545_), .C(_4307_), .Y(_4641_) );
	INVX1 INVX1_542 ( .A(_4404_), .Y(_4642_) );
	AOI22X1 AOI22X1_669 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_4315_), .C(_4642_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_4643_) );
	INVX1 INVX1_543 ( .A(_4416_), .Y(_4644_) );
	AOI22X1 AOI22X1_670 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_4451_), .C(_4644_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_4645_) );
	NAND3X1 NAND3X1_209 ( .A(_4645_), .B(_4641_), .C(_4643_), .Y(_4646_) );
	AOI22X1 AOI22X1_671 ( .A(_4400_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_4550_), .Y(_4647_) );
	AOI22X1 AOI22X1_672 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_4349_), .C(_4322_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_4648_) );
	INVX1 INVX1_544 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_4649_) );
	NAND2X1 NAND2X1_875 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_4439_), .Y(_4650_) );
	OAI21X1 OAI21X1_142 ( .A(_4649_), .B(_4411_), .C(_4650_), .Y(_4651_) );
	INVX1 INVX1_545 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_4652_) );
	NAND2X1 NAND2X1_876 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_4365_), .Y(_4653_) );
	OAI21X1 OAI21X1_143 ( .A(_4652_), .B(_4368_), .C(_4653_), .Y(_4654_) );
	NOR2X1 NOR2X1_508 ( .A(_4651_), .B(_4654_), .Y(_4655_) );
	NAND3X1 NAND3X1_210 ( .A(_4647_), .B(_4648_), .C(_4655_), .Y(_4656_) );
	INVX1 INVX1_546 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_4657_) );
	NAND2X1 NAND2X1_877 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_4347_), .Y(_4658_) );
	OAI21X1 OAI21X1_144 ( .A(_4657_), .B(_4377_), .C(_4658_), .Y(_4659_) );
	INVX1 INVX1_547 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_4660_) );
	INVX1 INVX1_548 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_4661_) );
	OAI22X1 OAI22X1_115 ( .A(_4660_), .B(_4383_), .C(_4381_), .D(_4661_), .Y(_4662_) );
	NOR2X1 NOR2X1_509 ( .A(_4662_), .B(_4659_), .Y(_4663_) );
	AOI22X1 AOI22X1_673 ( .A(_4467_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_4440_), .Y(_4664_) );
	AND2X2 AND2X2_93 ( .A(_4339_), .B(_4361_), .Y(_4665_) );
	AOI22X1 AOI22X1_674 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_4665_), .C(_4569_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_4666_) );
	NAND3X1 NAND3X1_211 ( .A(_4664_), .B(_4666_), .C(_4663_), .Y(_4667_) );
	NOR3X1 NOR3X1_367 ( .A(_4667_), .B(_4646_), .C(_4656_), .Y(_4668_) );
	INVX1 INVX1_549 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_4669_) );
	NOR3X1 NOR3X1_368 ( .A(_4669_), .B(_4334_), .C(_4333_), .Y(_4670_) );
	AND2X2 AND2X2_94 ( .A(_4355_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_4671_) );
	AND2X2 AND2X2_95 ( .A(_4475_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_4672_) );
	NOR3X1 NOR3X1_369 ( .A(_4672_), .B(_4671_), .C(_4670_), .Y(_4673_) );
	INVX1 INVX1_550 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_4674_) );
	INVX1 INVX1_551 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_4675_) );
	OAI22X1 OAI22X1_116 ( .A(_4675_), .B(_4410_), .C(_4360_), .D(_4674_), .Y(_4676_) );
	INVX1 INVX1_552 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_4677_) );
	INVX1 INVX1_553 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_4678_) );
	NAND2X1 NAND2X1_878 ( .A(_4351_), .B(_4352_), .Y(_4679_) );
	OAI22X1 OAI22X1_117 ( .A(_4679_), .B(_4678_), .C(_4677_), .D(_4330_), .Y(_4680_) );
	NOR2X1 NOR2X1_510 ( .A(_4676_), .B(_4680_), .Y(_4681_) );
	INVX1 INVX1_554 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_4682_) );
	NOR3X1 NOR3X1_370 ( .A(_4311_), .B(_4328_), .C(_4319_), .Y(_4683_) );
	NAND2X1 NAND2X1_879 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_4683_), .Y(_4684_) );
	OAI21X1 OAI21X1_145 ( .A(_4340_), .B(_4682_), .C(_4684_), .Y(_4685_) );
	INVX1 INVX1_555 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_4686_) );
	INVX1 INVX1_556 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_4687_) );
	OAI22X1 OAI22X1_118 ( .A(_4427_), .B(_4687_), .C(_4686_), .D(_4428_), .Y(_4688_) );
	NOR2X1 NOR2X1_511 ( .A(_4685_), .B(_4688_), .Y(_4689_) );
	NAND3X1 NAND3X1_212 ( .A(_4673_), .B(_4689_), .C(_4681_), .Y(_4690_) );
	AOI22X1 AOI22X1_675 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_4432_), .C(_4433_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_4691_) );
	AOI22X1 AOI22X1_676 ( .A(_4435_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_4436_), .Y(_4692_) );
	NAND2X1 NAND2X1_880 ( .A(_4691_), .B(_4692_), .Y(_4693_) );
	AOI22X1 AOI22X1_677 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_4443_), .C(_4442_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_4694_) );
	AOI22X1 AOI22X1_678 ( .A(_4386_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_4393_), .Y(_4695_) );
	NAND2X1 NAND2X1_881 ( .A(_4694_), .B(_4695_), .Y(_4696_) );
	NOR2X1 NOR2X1_512 ( .A(_4693_), .B(_4696_), .Y(_4697_) );
	AOI22X1 AOI22X1_679 ( .A(_4447_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_4448_), .Y(_4698_) );
	AOI22X1 AOI22X1_680 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_4474_), .C(_4450_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_4699_) );
	NAND2X1 NAND2X1_882 ( .A(_4699_), .B(_4698_), .Y(_4700_) );
	AOI22X1 AOI22X1_681 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_4454_), .C(_4455_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_4701_) );
	AOI22X1 AOI22X1_682 ( .A(_4457_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_4458_), .Y(_4702_) );
	NAND2X1 NAND2X1_883 ( .A(_4702_), .B(_4701_), .Y(_4703_) );
	NOR2X1 NOR2X1_513 ( .A(_4700_), .B(_4703_), .Y(_4704_) );
	NAND2X1 NAND2X1_884 ( .A(_4704_), .B(_4697_), .Y(_4705_) );
	AOI22X1 AOI22X1_683 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_4464_), .C(_4463_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_4706_) );
	AOI22X1 AOI22X1_684 ( .A(_4388_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_4466_), .Y(_4707_) );
	NAND2X1 NAND2X1_885 ( .A(_4706_), .B(_4707_), .Y(_4708_) );
	AOI22X1 AOI22X1_685 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_4472_), .C(_4470_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_4709_) );
	AOI22X1 AOI22X1_686 ( .A(_4402_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_4420_), .Y(_4710_) );
	NAND2X1 NAND2X1_886 ( .A(_4710_), .B(_4709_), .Y(_4711_) );
	NOR2X1 NOR2X1_514 ( .A(_4711_), .B(_4708_), .Y(_4712_) );
	AOI22X1 AOI22X1_687 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_4479_), .C(_4480_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_4713_) );
	NAND2X1 NAND2X1_887 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_4482_), .Y(_4714_) );
	NAND2X1 NAND2X1_888 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_4484_), .Y(_4715_) );
	NAND3X1 NAND3X1_213 ( .A(_4714_), .B(_4715_), .C(_4713_), .Y(_4716_) );
	AOI22X1 AOI22X1_688 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_4488_), .C(_4487_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_4717_) );
	AOI22X1 AOI22X1_689 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_4491_), .C(_4490_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_4718_) );
	NAND2X1 NAND2X1_889 ( .A(_4717_), .B(_4718_), .Y(_4719_) );
	NOR2X1 NOR2X1_515 ( .A(_4719_), .B(_4716_), .Y(_4720_) );
	NAND2X1 NAND2X1_890 ( .A(_4712_), .B(_4720_), .Y(_4721_) );
	NOR3X1 NOR3X1_371 ( .A(_4705_), .B(_4690_), .C(_4721_), .Y(_4722_) );
	AOI22X1 AOI22X1_690 ( .A(_4528_), .B(wData[42]), .C(wData[38]), .D(_4530_), .Y(_4723_) );
	AOI22X1 AOI22X1_691 ( .A(_4525_), .B(wData[46]), .C(_4532_), .D(wData[2]), .Y(_4724_) );
	NAND2X1 NAND2X1_891 ( .A(_4723_), .B(_4724_), .Y(_4725_) );
	AOI21X1 AOI21X1_102 ( .A(wData[34]), .B(_4518_), .C(_4725_), .Y(_4726_) );
	INVX1 INVX1_557 ( .A(wData[50]), .Y(_4727_) );
	AOI22X1 AOI22X1_692 ( .A(_4538_), .B(wData[10]), .C(wData[14]), .D(_4539_), .Y(_4728_) );
	OAI21X1 OAI21X1_146 ( .A(_4727_), .B(_4537_), .C(_4728_), .Y(_4729_) );
	AOI22X1 AOI22X1_693 ( .A(_4501_), .B(wData[22]), .C(wData[18]), .D(_4504_), .Y(_4730_) );
	NAND2X1 NAND2X1_892 ( .A(wData[26]), .B(_4508_), .Y(_4731_) );
	AOI22X1 AOI22X1_694 ( .A(_4514_), .B(wData[30]), .C(wData[6]), .D(_4512_), .Y(_4732_) );
	NAND3X1 NAND3X1_214 ( .A(_4731_), .B(_4732_), .C(_4730_), .Y(_4733_) );
	NOR2X1 NOR2X1_516 ( .A(_4729_), .B(_4733_), .Y(_4734_) );
	NAND2X1 NAND2X1_893 ( .A(wData[58]), .B(_4521_), .Y(_4735_) );
	NAND2X1 NAND2X1_894 ( .A(wData[54]), .B(_4522_), .Y(_4736_) );
	NAND2X1 NAND2X1_895 ( .A(_4735_), .B(_4736_), .Y(_4737_) );
	AOI21X1 AOI21X1_103 ( .A(wData[62]), .B(_4524_), .C(_4737_), .Y(_4738_) );
	NAND3X1 NAND3X1_215 ( .A(_4726_), .B(_4738_), .C(_4734_), .Y(_4739_) );
	NOR2X1 NOR2X1_517 ( .A(_4306_), .B(_4739_), .Y(_4740_) );
	AOI21X1 AOI21X1_104 ( .A(_4668_), .B(_4722_), .C(_4740_), .Y(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_2_) );
	AOI21X1 AOI21X1_105 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_4550_), .C(_4307_), .Y(_4741_) );
	AOI22X1 AOI22X1_695 ( .A(_4322_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_4642_), .Y(_4742_) );
	AOI22X1 AOI22X1_696 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_4644_), .C(_4400_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_4743_) );
	NAND3X1 NAND3X1_216 ( .A(_4743_), .B(_4741_), .C(_4742_), .Y(_4744_) );
	AOI22X1 AOI22X1_697 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_4349_), .C(_4347_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_4745_) );
	AOI22X1 AOI22X1_698 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_4420_), .C(_4545_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_4746_) );
	INVX1 INVX1_558 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_4747_) );
	INVX1 INVX1_559 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_4748_) );
	OAI22X1 OAI22X1_119 ( .A(_4747_), .B(_4362_), .C(_4411_), .D(_4748_), .Y(_4749_) );
	INVX1 INVX1_560 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_4750_) );
	NAND2X1 NAND2X1_896 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_4463_), .Y(_4751_) );
	OAI21X1 OAI21X1_147 ( .A(_4750_), .B(_4368_), .C(_4751_), .Y(_4752_) );
	NOR2X1 NOR2X1_518 ( .A(_4749_), .B(_4752_), .Y(_4753_) );
	NAND3X1 NAND3X1_217 ( .A(_4745_), .B(_4746_), .C(_4753_), .Y(_4754_) );
	AND2X2 AND2X2_96 ( .A(_4376_), .B(_4310_), .Y(_4755_) );
	AOI22X1 AOI22X1_699 ( .A(_4315_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_4755_), .Y(_4756_) );
	AND2X2 AND2X2_97 ( .A(_4374_), .B(_4339_), .Y(_4757_) );
	AND2X2 AND2X2_98 ( .A(_4382_), .B(_4339_), .Y(_4758_) );
	AOI22X1 AOI22X1_700 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_4758_), .C(_4757_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_4759_) );
	NAND2X1 NAND2X1_897 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_4467_), .Y(_4760_) );
	NAND2X1 NAND2X1_898 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_4440_), .Y(_4761_) );
	NAND2X1 NAND2X1_899 ( .A(_4760_), .B(_4761_), .Y(_4762_) );
	INVX1 INVX1_561 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_4763_) );
	NAND2X1 NAND2X1_900 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_4439_), .Y(_4764_) );
	OAI21X1 OAI21X1_148 ( .A(_4763_), .B(_4392_), .C(_4764_), .Y(_4765_) );
	NOR2X1 NOR2X1_519 ( .A(_4762_), .B(_4765_), .Y(_4766_) );
	NAND3X1 NAND3X1_218 ( .A(_4756_), .B(_4759_), .C(_4766_), .Y(_4767_) );
	NOR3X1 NOR3X1_372 ( .A(_4754_), .B(_4744_), .C(_4767_), .Y(_4768_) );
	INVX1 INVX1_562 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_4769_) );
	NAND2X1 NAND2X1_901 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_4355_), .Y(_4770_) );
	OAI21X1 OAI21X1_149 ( .A(_4360_), .B(_4769_), .C(_4770_), .Y(_4771_) );
	AOI21X1 AOI21X1_106 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_4335_), .C(_4771_), .Y(_4772_) );
	INVX1 INVX1_563 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_4773_) );
	INVX1 INVX1_564 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_4774_) );
	OAI22X1 OAI22X1_120 ( .A(_4679_), .B(_4774_), .C(_4773_), .D(_4330_), .Y(_4775_) );
	INVX1 INVX1_565 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_4776_) );
	NAND2X1 NAND2X1_902 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_4475_), .Y(_4777_) );
	OAI21X1 OAI21X1_150 ( .A(_4340_), .B(_4776_), .C(_4777_), .Y(_4778_) );
	NOR2X1 NOR2X1_520 ( .A(_4778_), .B(_4775_), .Y(_4779_) );
	INVX1 INVX1_566 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_4780_) );
	INVX1 INVX1_567 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_4781_) );
	OAI22X1 OAI22X1_121 ( .A(_4427_), .B(_4781_), .C(_4780_), .D(_4428_), .Y(_4782_) );
	INVX1 INVX1_568 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_4783_) );
	NAND2X1 NAND2X1_903 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_4474_), .Y(_4784_) );
	OAI21X1 OAI21X1_151 ( .A(_4783_), .B(_4410_), .C(_4784_), .Y(_4785_) );
	NOR2X1 NOR2X1_521 ( .A(_4785_), .B(_4782_), .Y(_4786_) );
	NAND3X1 NAND3X1_219 ( .A(_4772_), .B(_4786_), .C(_4779_), .Y(_4787_) );
	AOI22X1 AOI22X1_701 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_4432_), .C(_4433_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_4788_) );
	AOI22X1 AOI22X1_702 ( .A(_4435_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_4436_), .Y(_4789_) );
	NAND2X1 NAND2X1_904 ( .A(_4788_), .B(_4789_), .Y(_4790_) );
	AOI22X1 AOI22X1_703 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_4443_), .C(_4442_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_4791_) );
	AOI22X1 AOI22X1_704 ( .A(_4386_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_4393_), .Y(_4792_) );
	NAND2X1 NAND2X1_905 ( .A(_4791_), .B(_4792_), .Y(_4793_) );
	NOR2X1 NOR2X1_522 ( .A(_4790_), .B(_4793_), .Y(_4794_) );
	AOI22X1 AOI22X1_705 ( .A(_4447_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_4448_), .Y(_4795_) );
	AOI22X1 AOI22X1_706 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_4683_), .C(_4450_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_4796_) );
	NAND2X1 NAND2X1_906 ( .A(_4796_), .B(_4795_), .Y(_4797_) );
	AOI22X1 AOI22X1_707 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_4454_), .C(_4455_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_4798_) );
	AOI22X1 AOI22X1_708 ( .A(_4457_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_4458_), .Y(_4799_) );
	NAND2X1 NAND2X1_907 ( .A(_4799_), .B(_4798_), .Y(_4800_) );
	NOR2X1 NOR2X1_523 ( .A(_4797_), .B(_4800_), .Y(_4801_) );
	NAND2X1 NAND2X1_908 ( .A(_4801_), .B(_4794_), .Y(_4802_) );
	AOI22X1 AOI22X1_709 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_4464_), .C(_4365_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_4803_) );
	AOI22X1 AOI22X1_710 ( .A(_4388_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_4466_), .Y(_4804_) );
	NAND2X1 NAND2X1_909 ( .A(_4803_), .B(_4804_), .Y(_4805_) );
	AOI22X1 AOI22X1_711 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_4472_), .C(_4470_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_4806_) );
	AOI22X1 AOI22X1_712 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_4402_), .C(_4451_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_4807_) );
	NAND2X1 NAND2X1_910 ( .A(_4807_), .B(_4806_), .Y(_4808_) );
	NOR2X1 NOR2X1_524 ( .A(_4808_), .B(_4805_), .Y(_4809_) );
	AOI22X1 AOI22X1_713 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_4479_), .C(_4480_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_4810_) );
	NAND2X1 NAND2X1_911 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_4482_), .Y(_4811_) );
	NAND2X1 NAND2X1_912 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_4484_), .Y(_4812_) );
	NAND3X1 NAND3X1_220 ( .A(_4811_), .B(_4812_), .C(_4810_), .Y(_4813_) );
	AOI22X1 AOI22X1_714 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_4488_), .C(_4487_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_4814_) );
	AOI22X1 AOI22X1_715 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_4491_), .C(_4490_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_4815_) );
	NAND2X1 NAND2X1_913 ( .A(_4814_), .B(_4815_), .Y(_4816_) );
	NOR2X1 NOR2X1_525 ( .A(_4816_), .B(_4813_), .Y(_4817_) );
	NAND2X1 NAND2X1_914 ( .A(_4809_), .B(_4817_), .Y(_4818_) );
	NOR3X1 NOR3X1_373 ( .A(_4802_), .B(_4787_), .C(_4818_), .Y(_4819_) );
	NAND2X1 NAND2X1_915 ( .A(wData[59]), .B(_4521_), .Y(_4820_) );
	OAI21X1 OAI21X1_152 ( .A(_4305_), .B(wBusy_bF_buf0), .C(_4820_), .Y(_4821_) );
	NAND2X1 NAND2X1_916 ( .A(wData[7]), .B(_4512_), .Y(_4822_) );
	NAND2X1 NAND2X1_917 ( .A(wData[55]), .B(_4522_), .Y(_4823_) );
	AOI22X1 AOI22X1_716 ( .A(wData[63]), .B(_4524_), .C(_4514_), .D(wData[31]), .Y(_4824_) );
	NAND3X1 NAND3X1_221 ( .A(_4822_), .B(_4823_), .C(_4824_), .Y(_4825_) );
	OR2X2 OR2X2_50 ( .A(_4825_), .B(_4821_), .Y(_4826_) );
	INVX1 INVX1_569 ( .A(wData[51]), .Y(_4827_) );
	NAND2X1 NAND2X1_918 ( .A(wData[47]), .B(_4525_), .Y(_4828_) );
	OAI21X1 OAI21X1_153 ( .A(_4827_), .B(_4537_), .C(_4828_), .Y(_4829_) );
	AOI21X1 AOI21X1_107 ( .A(wData[3]), .B(_4532_), .C(_4829_), .Y(_4830_) );
	AOI22X1 AOI22X1_717 ( .A(_4538_), .B(wData[11]), .C(wData[15]), .D(_4539_), .Y(_4831_) );
	AOI22X1 AOI22X1_718 ( .A(_4501_), .B(wData[23]), .C(wData[27]), .D(_4508_), .Y(_4832_) );
	AND2X2 AND2X2_99 ( .A(_4831_), .B(_4832_), .Y(_4833_) );
	NAND2X1 NAND2X1_919 ( .A(wData[39]), .B(_4530_), .Y(_4834_) );
	NAND2X1 NAND2X1_920 ( .A(wData[43]), .B(_4528_), .Y(_4835_) );
	NAND2X1 NAND2X1_921 ( .A(_4834_), .B(_4835_), .Y(_4836_) );
	NAND2X1 NAND2X1_922 ( .A(wData[19]), .B(_4504_), .Y(_4837_) );
	NAND2X1 NAND2X1_923 ( .A(wData[35]), .B(_4518_), .Y(_4838_) );
	NAND2X1 NAND2X1_924 ( .A(_4837_), .B(_4838_), .Y(_4839_) );
	NOR2X1 NOR2X1_526 ( .A(_4836_), .B(_4839_), .Y(_4840_) );
	NAND3X1 NAND3X1_222 ( .A(_4833_), .B(_4830_), .C(_4840_), .Y(_4841_) );
	NOR2X1 NOR2X1_527 ( .A(_4826_), .B(_4841_), .Y(_4842_) );
	AOI21X1 AOI21X1_108 ( .A(_4768_), .B(_4819_), .C(_4842_), .Y(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_3_) );
	INVX1 INVX1_570 ( .A(wSelec[99]), .Y(_4843_) );
	NOR2X1 NOR2X1_528 ( .A(wBusy_bF_buf4), .B(_4843_), .Y(_4844_) );
	INVX1 INVX1_571 ( .A(_4844_), .Y(_4845_) );
	INVX1 INVX1_572 ( .A(wSelec[109]), .Y(_4846_) );
	NAND2X1 NAND2X1_925 ( .A(wSelec[108]), .B(_4846_), .Y(_4847_) );
	INVX2 INVX2_15 ( .A(_4847_), .Y(_4848_) );
	OR2X2 OR2X2_51 ( .A(wSelec[105]), .B(wSelec[104]), .Y(_4849_) );
	INVX1 INVX1_573 ( .A(wSelec[107]), .Y(_4850_) );
	NAND2X1 NAND2X1_926 ( .A(wSelec[106]), .B(_4850_), .Y(_4851_) );
	NOR2X1 NOR2X1_529 ( .A(_4849_), .B(_4851_), .Y(_4852_) );
	AND2X2 AND2X2_100 ( .A(_4852_), .B(_4848_), .Y(_4853_) );
	AOI21X1 AOI21X1_109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_4853_), .C(_4845_), .Y(_4854_) );
	INVX1 INVX1_574 ( .A(wSelec[105]), .Y(_4855_) );
	NAND2X1 NAND2X1_927 ( .A(wSelec[104]), .B(_4855_), .Y(_4856_) );
	OR2X2 OR2X2_52 ( .A(wSelec[106]), .B(wSelec[107]), .Y(_4857_) );
	NOR2X1 NOR2X1_530 ( .A(_4857_), .B(_4856_), .Y(_4858_) );
	NAND2X1 NAND2X1_928 ( .A(_4848_), .B(_4858_), .Y(_4859_) );
	INVX1 INVX1_575 ( .A(_4859_), .Y(_4860_) );
	INVX1 INVX1_576 ( .A(wSelec[104]), .Y(_4861_) );
	NAND2X1 NAND2X1_929 ( .A(wSelec[105]), .B(_4861_), .Y(_4862_) );
	INVX1 INVX1_577 ( .A(wSelec[106]), .Y(_4863_) );
	NAND2X1 NAND2X1_930 ( .A(wSelec[107]), .B(_4863_), .Y(_4864_) );
	NOR2X1 NOR2X1_531 ( .A(_4862_), .B(_4864_), .Y(_4865_) );
	NAND2X1 NAND2X1_931 ( .A(wSelec[108]), .B(wSelec[109]), .Y(_4866_) );
	INVX1 INVX1_578 ( .A(_4866_), .Y(_4867_) );
	NAND2X1 NAND2X1_932 ( .A(_4867_), .B(_4865_), .Y(_4868_) );
	INVX1 INVX1_579 ( .A(_4868_), .Y(_4869_) );
	AOI22X1 AOI22X1_719 ( .A(_4860_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_4869_), .Y(_4870_) );
	OR2X2 OR2X2_53 ( .A(_4856_), .B(_4857_), .Y(_4871_) );
	OR2X2 OR2X2_54 ( .A(wSelec[108]), .B(wSelec[109]), .Y(_4872_) );
	NOR2X1 NOR2X1_532 ( .A(_4872_), .B(_4871_), .Y(_4873_) );
	NOR2X1 NOR2X1_533 ( .A(_4851_), .B(_4856_), .Y(_4874_) );
	INVX1 INVX1_580 ( .A(wSelec[108]), .Y(_4875_) );
	NAND2X1 NAND2X1_933 ( .A(wSelec[109]), .B(_4875_), .Y(_4876_) );
	INVX2 INVX2_16 ( .A(_4876_), .Y(_4877_) );
	NAND2X1 NAND2X1_934 ( .A(_4877_), .B(_4874_), .Y(_4878_) );
	INVX1 INVX1_581 ( .A(_4878_), .Y(_4879_) );
	AOI22X1 AOI22X1_720 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_4873_), .C(_4879_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_4880_) );
	NAND3X1 NAND3X1_223 ( .A(_4854_), .B(_4880_), .C(_4870_), .Y(_4881_) );
	NOR2X1 NOR2X1_534 ( .A(wSelec[105]), .B(wSelec[104]), .Y(_4882_) );
	NOR2X1 NOR2X1_535 ( .A(wSelec[106]), .B(wSelec[107]), .Y(_4883_) );
	NAND2X1 NAND2X1_935 ( .A(_4882_), .B(_4883_), .Y(_4884_) );
	NOR2X1 NOR2X1_536 ( .A(_4847_), .B(_4884_), .Y(_4885_) );
	NAND2X1 NAND2X1_936 ( .A(wSelec[105]), .B(wSelec[104]), .Y(_4886_) );
	NOR3X1 NOR3X1_374 ( .A(_4857_), .B(_4886_), .C(_4847_), .Y(_4887_) );
	AOI22X1 AOI22X1_721 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_4887_), .C(_4885_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_4888_) );
	INVX1 INVX1_582 ( .A(_4872_), .Y(_4889_) );
	NOR2X1 NOR2X1_537 ( .A(_4857_), .B(_4862_), .Y(_4890_) );
	AND2X2 AND2X2_101 ( .A(_4890_), .B(_4889_), .Y(_4891_) );
	NAND2X1 NAND2X1_937 ( .A(wSelec[106]), .B(wSelec[107]), .Y(_4892_) );
	NOR3X1 NOR3X1_375 ( .A(_4866_), .B(_4886_), .C(_4892_), .Y(_4893_) );
	AOI22X1 AOI22X1_722 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_4893_), .C(_4891_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_4894_) );
	INVX1 INVX1_583 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_4895_) );
	INVX1 INVX1_584 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_4896_) );
	NOR2X1 NOR2X1_538 ( .A(_4856_), .B(_4864_), .Y(_4897_) );
	NAND2X1 NAND2X1_938 ( .A(_4867_), .B(_4897_), .Y(_4898_) );
	NOR2X1 NOR2X1_539 ( .A(_4886_), .B(_4892_), .Y(_4899_) );
	NAND2X1 NAND2X1_939 ( .A(_4899_), .B(_4877_), .Y(_4900_) );
	OAI22X1 OAI22X1_122 ( .A(_4895_), .B(_4900_), .C(_4898_), .D(_4896_), .Y(_4901_) );
	INVX1 INVX1_585 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_4902_) );
	NOR3X1 NOR3X1_376 ( .A(_4847_), .B(_4862_), .C(_4864_), .Y(_4903_) );
	NAND2X1 NAND2X1_940 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_4903_), .Y(_4904_) );
	NOR2X1 NOR2X1_540 ( .A(_4886_), .B(_4851_), .Y(_4905_) );
	NAND2X1 NAND2X1_941 ( .A(_4877_), .B(_4905_), .Y(_4906_) );
	OAI21X1 OAI21X1_154 ( .A(_4902_), .B(_4906_), .C(_4904_), .Y(_4907_) );
	NOR2X1 NOR2X1_541 ( .A(_4901_), .B(_4907_), .Y(_4908_) );
	NAND3X1 NAND3X1_224 ( .A(_4888_), .B(_4894_), .C(_4908_), .Y(_4909_) );
	INVX1 INVX1_586 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_4910_) );
	INVX1 INVX1_587 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_4911_) );
	NOR2X1 NOR2X1_542 ( .A(_4851_), .B(_4862_), .Y(_4912_) );
	NAND2X1 NAND2X1_942 ( .A(_4848_), .B(_4912_), .Y(_4913_) );
	NOR2X1 NOR2X1_543 ( .A(_4849_), .B(_4864_), .Y(_4914_) );
	NAND2X1 NAND2X1_943 ( .A(_4848_), .B(_4914_), .Y(_4915_) );
	OAI22X1 OAI22X1_123 ( .A(_4915_), .B(_4910_), .C(_4911_), .D(_4913_), .Y(_4916_) );
	INVX1 INVX1_588 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_4917_) );
	INVX1 INVX1_589 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_4918_) );
	NAND2X1 NAND2X1_944 ( .A(_4877_), .B(_4912_), .Y(_4919_) );
	NOR2X1 NOR2X1_544 ( .A(_4886_), .B(_4857_), .Y(_4920_) );
	NAND2X1 NAND2X1_945 ( .A(_4877_), .B(_4920_), .Y(_4921_) );
	OAI22X1 OAI22X1_124 ( .A(_4917_), .B(_4921_), .C(_4919_), .D(_4918_), .Y(_4922_) );
	NOR2X1 NOR2X1_545 ( .A(_4922_), .B(_4916_), .Y(_4923_) );
	NOR3X1 NOR3X1_377 ( .A(_4856_), .B(_4892_), .C(_4876_), .Y(_4924_) );
	NAND2X1 NAND2X1_946 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_4924_), .Y(_4925_) );
	NOR3X1 NOR3X1_378 ( .A(_4864_), .B(_4886_), .C(_4876_), .Y(_4926_) );
	NAND2X1 NAND2X1_947 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_4926_), .Y(_4927_) );
	NAND2X1 NAND2X1_948 ( .A(_4925_), .B(_4927_), .Y(_4928_) );
	INVX1 INVX1_590 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_4929_) );
	NAND2X1 NAND2X1_949 ( .A(_4867_), .B(_4852_), .Y(_4930_) );
	NOR3X1 NOR3X1_379 ( .A(_4862_), .B(_4864_), .C(_4876_), .Y(_4931_) );
	NAND2X1 NAND2X1_950 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_4931_), .Y(_4932_) );
	OAI21X1 OAI21X1_155 ( .A(_4929_), .B(_4930_), .C(_4932_), .Y(_4933_) );
	NOR2X1 NOR2X1_546 ( .A(_4928_), .B(_4933_), .Y(_4934_) );
	NAND2X1 NAND2X1_951 ( .A(_4923_), .B(_4934_), .Y(_4935_) );
	NOR3X1 NOR3X1_380 ( .A(_4881_), .B(_4935_), .C(_4909_), .Y(_4936_) );
	NAND2X1 NAND2X1_952 ( .A(_4848_), .B(_4905_), .Y(_4937_) );
	INVX1 INVX1_591 ( .A(_4937_), .Y(_4938_) );
	INVX1 INVX1_592 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_4939_) );
	NOR3X1 NOR3X1_381 ( .A(_4849_), .B(_4872_), .C(_4851_), .Y(_4940_) );
	NAND2X1 NAND2X1_953 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_4940_), .Y(_4941_) );
	NAND2X1 NAND2X1_954 ( .A(_4889_), .B(_4912_), .Y(_4942_) );
	OAI21X1 OAI21X1_156 ( .A(_4942_), .B(_4939_), .C(_4941_), .Y(_4943_) );
	AOI21X1 AOI21X1_110 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_4938_), .C(_4943_), .Y(_4944_) );
	INVX1 INVX1_593 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_4945_) );
	INVX1 INVX1_594 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_4946_) );
	NOR2X1 NOR2X1_547 ( .A(_4892_), .B(_4849_), .Y(_4947_) );
	NAND2X1 NAND2X1_955 ( .A(_4848_), .B(_4947_), .Y(_4948_) );
	NAND2X1 NAND2X1_956 ( .A(_4889_), .B(_4874_), .Y(_4949_) );
	OAI22X1 OAI22X1_125 ( .A(_4946_), .B(_4948_), .C(_4949_), .D(_4945_), .Y(_4950_) );
	INVX1 INVX1_595 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_4951_) );
	INVX1 INVX1_596 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_4952_) );
	NAND2X1 NAND2X1_957 ( .A(_4848_), .B(_4874_), .Y(_4953_) );
	NAND2X1 NAND2X1_958 ( .A(_4889_), .B(_4920_), .Y(_4954_) );
	OAI22X1 OAI22X1_126 ( .A(_4951_), .B(_4954_), .C(_4953_), .D(_4952_), .Y(_4955_) );
	NOR2X1 NOR2X1_548 ( .A(_4950_), .B(_4955_), .Y(_4956_) );
	INVX1 INVX1_597 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_4957_) );
	NOR3X1 NOR3X1_382 ( .A(_4872_), .B(_4886_), .C(_4851_), .Y(_4958_) );
	NAND2X1 NAND2X1_959 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_4958_), .Y(_4959_) );
	OR2X2 OR2X2_55 ( .A(_4884_), .B(_4866_), .Y(_4960_) );
	OAI21X1 OAI21X1_157 ( .A(_4957_), .B(_4960_), .C(_4959_), .Y(_4961_) );
	INVX1 INVX1_598 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_4962_) );
	INVX1 INVX1_599 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_4963_) );
	NOR2X1 NOR2X1_549 ( .A(_4892_), .B(_4862_), .Y(_4964_) );
	NAND2X1 NAND2X1_960 ( .A(_4848_), .B(_4964_), .Y(_4965_) );
	NAND2X1 NAND2X1_961 ( .A(_4867_), .B(_4858_), .Y(_4966_) );
	OAI22X1 OAI22X1_127 ( .A(_4965_), .B(_4963_), .C(_4962_), .D(_4966_), .Y(_4967_) );
	NOR2X1 NOR2X1_550 ( .A(_4961_), .B(_4967_), .Y(_4968_) );
	NAND3X1 NAND3X1_225 ( .A(_4944_), .B(_4968_), .C(_4956_), .Y(_4969_) );
	NOR3X1 NOR3X1_383 ( .A(_4849_), .B(_4857_), .C(_4872_), .Y(_4970_) );
	NOR3X1 NOR3X1_384 ( .A(_4866_), .B(_4892_), .C(_4856_), .Y(_4971_) );
	AOI22X1 AOI22X1_723 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_4970_), .C(_4971_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_4972_) );
	NOR3X1 NOR3X1_385 ( .A(_4866_), .B(_4892_), .C(_4862_), .Y(_4973_) );
	NOR3X1 NOR3X1_386 ( .A(_4866_), .B(_4886_), .C(_4864_), .Y(_4974_) );
	AOI22X1 AOI22X1_724 ( .A(_4973_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_4974_), .Y(_4975_) );
	NAND2X1 NAND2X1_962 ( .A(_4972_), .B(_4975_), .Y(_4976_) );
	NOR3X1 NOR3X1_387 ( .A(_4864_), .B(_4849_), .C(_4876_), .Y(_4977_) );
	NOR3X1 NOR3X1_388 ( .A(_4856_), .B(_4864_), .C(_4876_), .Y(_4978_) );
	AOI22X1 AOI22X1_725 ( .A(_4977_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_4978_), .Y(_4979_) );
	NOR3X1 NOR3X1_389 ( .A(_4847_), .B(_4892_), .C(_4856_), .Y(_4980_) );
	NOR3X1 NOR3X1_390 ( .A(_4886_), .B(_4892_), .C(_4847_), .Y(_4981_) );
	AOI22X1 AOI22X1_726 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_4981_), .C(_4980_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_4982_) );
	NAND2X1 NAND2X1_963 ( .A(_4982_), .B(_4979_), .Y(_4983_) );
	NOR2X1 NOR2X1_551 ( .A(_4976_), .B(_4983_), .Y(_4984_) );
	NOR3X1 NOR3X1_391 ( .A(_4872_), .B(_4892_), .C(_4856_), .Y(_4985_) );
	NOR3X1 NOR3X1_392 ( .A(_4872_), .B(_4892_), .C(_4862_), .Y(_4986_) );
	AOI22X1 AOI22X1_727 ( .A(_4985_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_4986_), .Y(_4987_) );
	NOR3X1 NOR3X1_393 ( .A(_4872_), .B(_4886_), .C(_4864_), .Y(_4988_) );
	NOR3X1 NOR3X1_394 ( .A(_4847_), .B(_4857_), .C(_4862_), .Y(_4989_) );
	AOI22X1 AOI22X1_728 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_4988_), .C(_4989_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_4990_) );
	NAND2X1 NAND2X1_964 ( .A(_4987_), .B(_4990_), .Y(_4991_) );
	NOR3X1 NOR3X1_395 ( .A(_4886_), .B(_4892_), .C(_4872_), .Y(_4992_) );
	NOR3X1 NOR3X1_396 ( .A(_4862_), .B(_4857_), .C(_4876_), .Y(_4993_) );
	AOI22X1 AOI22X1_729 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_4992_), .C(_4993_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_4994_) );
	NOR3X1 NOR3X1_397 ( .A(_4849_), .B(_4857_), .C(_4876_), .Y(_4995_) );
	NOR3X1 NOR3X1_398 ( .A(_4849_), .B(_4892_), .C(_4876_), .Y(_4996_) );
	AOI22X1 AOI22X1_730 ( .A(_4995_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_4996_), .Y(_4997_) );
	NAND2X1 NAND2X1_965 ( .A(_4997_), .B(_4994_), .Y(_4998_) );
	NOR2X1 NOR2X1_552 ( .A(_4991_), .B(_4998_), .Y(_4999_) );
	NAND2X1 NAND2X1_966 ( .A(_4999_), .B(_4984_), .Y(_5000_) );
	NOR3X1 NOR3X1_399 ( .A(_4847_), .B(_4886_), .C(_4864_), .Y(_5001_) );
	NOR3X1 NOR3X1_400 ( .A(_4857_), .B(_4866_), .C(_4862_), .Y(_5002_) );
	AOI22X1 AOI22X1_731 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_5002_), .C(_5001_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_5003_) );
	NOR3X1 NOR3X1_401 ( .A(_4851_), .B(_4849_), .C(_4876_), .Y(_5004_) );
	NOR3X1 NOR3X1_402 ( .A(_4862_), .B(_4892_), .C(_4876_), .Y(_5005_) );
	AOI22X1 AOI22X1_732 ( .A(_5004_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_5005_), .Y(_5006_) );
	NAND2X1 NAND2X1_967 ( .A(_5003_), .B(_5006_), .Y(_5007_) );
	NOR3X1 NOR3X1_403 ( .A(_4847_), .B(_4856_), .C(_4864_), .Y(_5008_) );
	NAND2X1 NAND2X1_968 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_5008_), .Y(_5009_) );
	NOR3X1 NOR3X1_404 ( .A(_4866_), .B(_4886_), .C(_4851_), .Y(_5010_) );
	NAND2X1 NAND2X1_969 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_5010_), .Y(_5011_) );
	NOR3X1 NOR3X1_405 ( .A(_4849_), .B(_4892_), .C(_4872_), .Y(_5012_) );
	NOR3X1 NOR3X1_406 ( .A(_4849_), .B(_4866_), .C(_4864_), .Y(_5013_) );
	AOI22X1 AOI22X1_733 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_5012_), .C(_5013_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_5014_) );
	NAND3X1 NAND3X1_226 ( .A(_5009_), .B(_5011_), .C(_5014_), .Y(_5015_) );
	NOR2X1 NOR2X1_553 ( .A(_5015_), .B(_5007_), .Y(_5016_) );
	NOR3X1 NOR3X1_407 ( .A(_4849_), .B(_4872_), .C(_4864_), .Y(_5017_) );
	NOR3X1 NOR3X1_408 ( .A(_4851_), .B(_4866_), .C(_4856_), .Y(_5018_) );
	AOI22X1 AOI22X1_734 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_5017_), .C(_5018_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_5019_) );
	NOR3X1 NOR3X1_409 ( .A(_4851_), .B(_4866_), .C(_4862_), .Y(_5020_) );
	NAND2X1 NAND2X1_970 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_5020_), .Y(_5021_) );
	NOR3X1 NOR3X1_410 ( .A(_4856_), .B(_4857_), .C(_4876_), .Y(_5022_) );
	NAND2X1 NAND2X1_971 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_5022_), .Y(_5023_) );
	NAND3X1 NAND3X1_227 ( .A(_5021_), .B(_5023_), .C(_5019_), .Y(_5024_) );
	NOR3X1 NOR3X1_411 ( .A(_4856_), .B(_4872_), .C(_4864_), .Y(_5025_) );
	NOR3X1 NOR3X1_412 ( .A(_4866_), .B(_4892_), .C(_4849_), .Y(_5026_) );
	AOI22X1 AOI22X1_735 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_5026_), .C(_5025_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_5027_) );
	NOR3X1 NOR3X1_413 ( .A(_4862_), .B(_4872_), .C(_4864_), .Y(_5028_) );
	NOR3X1 NOR3X1_414 ( .A(_4866_), .B(_4886_), .C(_4857_), .Y(_5029_) );
	AOI22X1 AOI22X1_736 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_5029_), .C(_5028_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_5030_) );
	NAND2X1 NAND2X1_972 ( .A(_5027_), .B(_5030_), .Y(_5031_) );
	NOR2X1 NOR2X1_554 ( .A(_5031_), .B(_5024_), .Y(_5032_) );
	NAND2X1 NAND2X1_973 ( .A(_5016_), .B(_5032_), .Y(_5033_) );
	NOR3X1 NOR3X1_415 ( .A(_5000_), .B(_4969_), .C(_5033_), .Y(_5034_) );
	INVX1 INVX1_600 ( .A(wSelec[101]), .Y(_5035_) );
	NAND2X1 NAND2X1_974 ( .A(wSelec[100]), .B(_5035_), .Y(_5036_) );
	INVX1 INVX1_601 ( .A(wSelec[103]), .Y(_5037_) );
	NAND2X1 NAND2X1_975 ( .A(wSelec[102]), .B(_5037_), .Y(_5038_) );
	NOR2X1 NOR2X1_555 ( .A(_5036_), .B(_5038_), .Y(_5039_) );
	NOR2X1 NOR2X1_556 ( .A(wSelec[101]), .B(wSelec[100]), .Y(_5040_) );
	INVX1 INVX1_602 ( .A(_5040_), .Y(_5041_) );
	NOR2X1 NOR2X1_557 ( .A(_5038_), .B(_5041_), .Y(_5042_) );
	AOI22X1 AOI22X1_737 ( .A(wData[20]), .B(_5039_), .C(_5042_), .D(wData[16]), .Y(_5043_) );
	INVX1 INVX1_603 ( .A(wSelec[100]), .Y(_5044_) );
	NAND2X1 NAND2X1_976 ( .A(wSelec[101]), .B(_5044_), .Y(_5045_) );
	NOR2X1 NOR2X1_558 ( .A(_5045_), .B(_5038_), .Y(_5046_) );
	NAND2X1 NAND2X1_977 ( .A(wData[24]), .B(_5046_), .Y(_5047_) );
	INVX1 INVX1_604 ( .A(wSelec[102]), .Y(_5048_) );
	NAND2X1 NAND2X1_978 ( .A(_5048_), .B(_5037_), .Y(_5049_) );
	NOR2X1 NOR2X1_559 ( .A(_5036_), .B(_5049_), .Y(_5050_) );
	NAND2X1 NAND2X1_979 ( .A(wSelec[101]), .B(wSelec[100]), .Y(_5051_) );
	NOR2X1 NOR2X1_560 ( .A(_5051_), .B(_5038_), .Y(_5052_) );
	AOI22X1 AOI22X1_738 ( .A(_5052_), .B(wData[28]), .C(wData[4]), .D(_5050_), .Y(_5053_) );
	NAND3X1 NAND3X1_228 ( .A(_5047_), .B(_5053_), .C(_5043_), .Y(_5054_) );
	NAND2X1 NAND2X1_980 ( .A(wSelec[103]), .B(_5048_), .Y(_5055_) );
	NOR2X1 NOR2X1_561 ( .A(_5055_), .B(_5041_), .Y(_5056_) );
	NAND2X1 NAND2X1_981 ( .A(wData[32]), .B(_5056_), .Y(_5057_) );
	NAND2X1 NAND2X1_982 ( .A(wSelec[102]), .B(wSelec[103]), .Y(_5058_) );
	NOR2X1 NOR2X1_562 ( .A(_5058_), .B(_5045_), .Y(_5059_) );
	NOR2X1 NOR2X1_563 ( .A(_5058_), .B(_5036_), .Y(_5060_) );
	AOI22X1 AOI22X1_739 ( .A(_5059_), .B(wData[56]), .C(wData[52]), .D(_5060_), .Y(_5061_) );
	NOR2X1 NOR2X1_564 ( .A(_5051_), .B(_5058_), .Y(_5062_) );
	NOR2X1 NOR2X1_565 ( .A(_5051_), .B(_5055_), .Y(_5063_) );
	AOI22X1 AOI22X1_740 ( .A(wData[60]), .B(_5062_), .C(_5063_), .D(wData[44]), .Y(_5064_) );
	NAND3X1 NAND3X1_229 ( .A(_5057_), .B(_5064_), .C(_5061_), .Y(_5065_) );
	NOR2X1 NOR2X1_566 ( .A(_5045_), .B(_5055_), .Y(_5066_) );
	NAND2X1 NAND2X1_983 ( .A(wData[40]), .B(_5066_), .Y(_5067_) );
	NOR2X1 NOR2X1_567 ( .A(_5055_), .B(_5036_), .Y(_5068_) );
	NAND2X1 NAND2X1_984 ( .A(wData[36]), .B(_5068_), .Y(_5069_) );
	NOR2X1 NOR2X1_568 ( .A(_5049_), .B(_5041_), .Y(_5070_) );
	NAND2X1 NAND2X1_985 ( .A(wData[0]), .B(_5070_), .Y(_5071_) );
	NAND3X1 NAND3X1_230 ( .A(_5067_), .B(_5069_), .C(_5071_), .Y(_5072_) );
	INVX1 INVX1_605 ( .A(wData[48]), .Y(_5073_) );
	NOR2X1 NOR2X1_569 ( .A(_5048_), .B(_5037_), .Y(_5074_) );
	NAND2X1 NAND2X1_986 ( .A(_5040_), .B(_5074_), .Y(_5075_) );
	NOR2X1 NOR2X1_570 ( .A(_5045_), .B(_5049_), .Y(_5076_) );
	NOR2X1 NOR2X1_571 ( .A(_5051_), .B(_5049_), .Y(_5077_) );
	AOI22X1 AOI22X1_741 ( .A(_5076_), .B(wData[8]), .C(wData[12]), .D(_5077_), .Y(_5078_) );
	OAI21X1 OAI21X1_158 ( .A(_5073_), .B(_5075_), .C(_5078_), .Y(_5079_) );
	OR2X2 OR2X2_56 ( .A(_5079_), .B(_5072_), .Y(_5080_) );
	NOR3X1 NOR3X1_416 ( .A(_5054_), .B(_5065_), .C(_5080_), .Y(_5081_) );
	AND2X2 AND2X2_102 ( .A(_5081_), .B(_4845_), .Y(_5082_) );
	AOI21X1 AOI21X1_111 ( .A(_4936_), .B(_5034_), .C(_5082_), .Y(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_0_) );
	INVX1 INVX1_606 ( .A(_4953_), .Y(_5083_) );
	AOI21X1 AOI21X1_112 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_5083_), .C(_4845_), .Y(_5084_) );
	AOI22X1 AOI22X1_742 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_4853_), .C(_4869_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_5085_) );
	AOI22X1 AOI22X1_743 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_4873_), .C(_4879_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_5086_) );
	NAND3X1 NAND3X1_231 ( .A(_5084_), .B(_5085_), .C(_5086_), .Y(_5087_) );
	INVX1 INVX1_607 ( .A(_4913_), .Y(_5088_) );
	AOI22X1 AOI22X1_744 ( .A(_4938_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_5088_), .Y(_5089_) );
	AOI22X1 AOI22X1_745 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_5012_), .C(_4891_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_5090_) );
	INVX1 INVX1_608 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_5091_) );
	INVX1 INVX1_609 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_5092_) );
	OAI22X1 OAI22X1_128 ( .A(_5091_), .B(_4900_), .C(_4898_), .D(_5092_), .Y(_5093_) );
	INVX1 INVX1_610 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_5094_) );
	NAND2X1 NAND2X1_987 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_5001_), .Y(_5095_) );
	OAI21X1 OAI21X1_159 ( .A(_5094_), .B(_4906_), .C(_5095_), .Y(_5096_) );
	NOR2X1 NOR2X1_572 ( .A(_5093_), .B(_5096_), .Y(_5097_) );
	NAND3X1 NAND3X1_232 ( .A(_5089_), .B(_5090_), .C(_5097_), .Y(_5098_) );
	INVX1 INVX1_611 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_5099_) );
	NAND2X1 NAND2X1_988 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_4885_), .Y(_5100_) );
	OAI21X1 OAI21X1_160 ( .A(_5099_), .B(_4915_), .C(_5100_), .Y(_5101_) );
	INVX1 INVX1_612 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_5102_) );
	INVX1 INVX1_613 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_5103_) );
	OAI22X1 OAI22X1_129 ( .A(_5102_), .B(_4921_), .C(_4919_), .D(_5103_), .Y(_5104_) );
	NOR2X1 NOR2X1_573 ( .A(_5104_), .B(_5101_), .Y(_5105_) );
	AOI22X1 AOI22X1_746 ( .A(_5005_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_4978_), .Y(_5106_) );
	AND2X2 AND2X2_103 ( .A(_4852_), .B(_4867_), .Y(_5107_) );
	AOI22X1 AOI22X1_747 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_4977_), .C(_5107_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_5108_) );
	NAND3X1 NAND3X1_233 ( .A(_5106_), .B(_5108_), .C(_5105_), .Y(_5109_) );
	NOR3X1 NOR3X1_417 ( .A(_5109_), .B(_5087_), .C(_5098_), .Y(_5110_) );
	INVX1 INVX1_614 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_5111_) );
	NAND2X1 NAND2X1_989 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_4940_), .Y(_5112_) );
	OAI21X1 OAI21X1_161 ( .A(_4942_), .B(_5111_), .C(_5112_), .Y(_5113_) );
	AOI21X1 AOI21X1_113 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_4989_), .C(_5113_), .Y(_5114_) );
	INVX1 INVX1_615 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_5115_) );
	INVX1 INVX1_616 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_5116_) );
	OAI22X1 OAI22X1_130 ( .A(_5116_), .B(_4948_), .C(_4949_), .D(_5115_), .Y(_5117_) );
	INVX1 INVX1_617 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_5118_) );
	NAND2X1 NAND2X1_990 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_4958_), .Y(_5119_) );
	OAI21X1 OAI21X1_162 ( .A(_4859_), .B(_5118_), .C(_5119_), .Y(_5120_) );
	NOR2X1 NOR2X1_574 ( .A(_5120_), .B(_5117_), .Y(_5121_) );
	INVX1 INVX1_618 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_5122_) );
	INVX1 INVX1_619 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_5123_) );
	OAI22X1 OAI22X1_131 ( .A(_4954_), .B(_5123_), .C(_4960_), .D(_5122_), .Y(_5124_) );
	INVX1 INVX1_620 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_5125_) );
	NOR2X1 NOR2X1_575 ( .A(_5125_), .B(_4965_), .Y(_5126_) );
	INVX1 INVX1_621 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_5127_) );
	NOR2X1 NOR2X1_576 ( .A(_5127_), .B(_4966_), .Y(_5128_) );
	NOR3X1 NOR3X1_418 ( .A(_5126_), .B(_5124_), .C(_5128_), .Y(_5129_) );
	NAND3X1 NAND3X1_234 ( .A(_5121_), .B(_5114_), .C(_5129_), .Y(_5130_) );
	AOI22X1 AOI22X1_748 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_4970_), .C(_4971_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_5131_) );
	AOI22X1 AOI22X1_749 ( .A(_4973_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_4974_), .Y(_5132_) );
	NAND2X1 NAND2X1_991 ( .A(_5131_), .B(_5132_), .Y(_5133_) );
	AOI22X1 AOI22X1_750 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_4981_), .C(_4980_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_5134_) );
	AOI22X1 AOI22X1_751 ( .A(_4924_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_4931_), .Y(_5135_) );
	NAND2X1 NAND2X1_992 ( .A(_5134_), .B(_5135_), .Y(_5136_) );
	NOR2X1 NOR2X1_577 ( .A(_5133_), .B(_5136_), .Y(_5137_) );
	AOI22X1 AOI22X1_752 ( .A(_4985_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_4986_), .Y(_5138_) );
	AOI22X1 AOI22X1_753 ( .A(_4887_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_4988_), .Y(_5139_) );
	NAND2X1 NAND2X1_993 ( .A(_5138_), .B(_5139_), .Y(_5140_) );
	AOI22X1 AOI22X1_754 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_4992_), .C(_4993_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_5141_) );
	AOI22X1 AOI22X1_755 ( .A(_4995_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_4996_), .Y(_5142_) );
	NAND2X1 NAND2X1_994 ( .A(_5142_), .B(_5141_), .Y(_5143_) );
	NOR2X1 NOR2X1_578 ( .A(_5140_), .B(_5143_), .Y(_5144_) );
	NAND2X1 NAND2X1_995 ( .A(_5144_), .B(_5137_), .Y(_5145_) );
	AOI22X1 AOI22X1_756 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_5002_), .C(_4903_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_5146_) );
	AOI22X1 AOI22X1_757 ( .A(_4926_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_5004_), .Y(_5147_) );
	NAND2X1 NAND2X1_996 ( .A(_5146_), .B(_5147_), .Y(_5148_) );
	AOI22X1 AOI22X1_758 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_4893_), .C(_5013_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_5149_) );
	NAND2X1 NAND2X1_997 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_5008_), .Y(_5150_) );
	NAND2X1 NAND2X1_998 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_5010_), .Y(_5151_) );
	NAND3X1 NAND3X1_235 ( .A(_5150_), .B(_5151_), .C(_5149_), .Y(_5152_) );
	NOR2X1 NOR2X1_579 ( .A(_5152_), .B(_5148_), .Y(_5153_) );
	AOI22X1 AOI22X1_759 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_5017_), .C(_5018_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_5154_) );
	NAND2X1 NAND2X1_999 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_5020_), .Y(_5155_) );
	NAND2X1 NAND2X1_1000 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_5022_), .Y(_5156_) );
	NAND3X1 NAND3X1_236 ( .A(_5155_), .B(_5156_), .C(_5154_), .Y(_5157_) );
	AOI22X1 AOI22X1_760 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_5026_), .C(_5025_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_5158_) );
	AOI22X1 AOI22X1_761 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_5029_), .C(_5028_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_5159_) );
	NAND2X1 NAND2X1_1001 ( .A(_5158_), .B(_5159_), .Y(_5160_) );
	NOR2X1 NOR2X1_580 ( .A(_5160_), .B(_5157_), .Y(_5161_) );
	NAND2X1 NAND2X1_1002 ( .A(_5153_), .B(_5161_), .Y(_5162_) );
	NOR3X1 NOR3X1_419 ( .A(_5145_), .B(_5130_), .C(_5162_), .Y(_5163_) );
	AOI21X1 AOI21X1_114 ( .A(wData[21]), .B(_5039_), .C(_4844_), .Y(_5164_) );
	AOI22X1 AOI22X1_762 ( .A(_5042_), .B(wData[17]), .C(wData[1]), .D(_5070_), .Y(_5165_) );
	AOI22X1 AOI22X1_763 ( .A(_5063_), .B(wData[45]), .C(wData[25]), .D(_5046_), .Y(_5166_) );
	NAND3X1 NAND3X1_237 ( .A(_5164_), .B(_5166_), .C(_5165_), .Y(_5167_) );
	NAND3X1 NAND3X1_238 ( .A(wData[49]), .B(_5040_), .C(_5074_), .Y(_5168_) );
	AOI22X1 AOI22X1_764 ( .A(wData[61]), .B(_5062_), .C(_5050_), .D(wData[5]), .Y(_5169_) );
	AND2X2 AND2X2_104 ( .A(_5169_), .B(_5168_), .Y(_5170_) );
	AOI22X1 AOI22X1_765 ( .A(_5059_), .B(wData[57]), .C(wData[41]), .D(_5066_), .Y(_5171_) );
	AOI22X1 AOI22X1_766 ( .A(wData[53]), .B(_5060_), .C(_5056_), .D(wData[33]), .Y(_5172_) );
	AND2X2 AND2X2_105 ( .A(_5172_), .B(_5171_), .Y(_5173_) );
	AOI22X1 AOI22X1_767 ( .A(_5076_), .B(wData[9]), .C(wData[13]), .D(_5077_), .Y(_5174_) );
	AOI22X1 AOI22X1_768 ( .A(_5052_), .B(wData[29]), .C(wData[37]), .D(_5068_), .Y(_5175_) );
	AND2X2 AND2X2_106 ( .A(_5174_), .B(_5175_), .Y(_5176_) );
	NAND3X1 NAND3X1_239 ( .A(_5170_), .B(_5176_), .C(_5173_), .Y(_5177_) );
	NOR2X1 NOR2X1_581 ( .A(_5167_), .B(_5177_), .Y(_5178_) );
	AOI21X1 AOI21X1_115 ( .A(_5110_), .B(_5163_), .C(_5178_), .Y(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_1_) );
	AOI21X1 AOI21X1_116 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_5083_), .C(_4845_), .Y(_5179_) );
	INVX1 INVX1_622 ( .A(_4942_), .Y(_5180_) );
	AOI22X1 AOI22X1_769 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_4853_), .C(_5180_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_5181_) );
	INVX1 INVX1_623 ( .A(_4954_), .Y(_5182_) );
	AOI22X1 AOI22X1_770 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_4989_), .C(_5182_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_5183_) );
	NAND3X1 NAND3X1_240 ( .A(_5183_), .B(_5179_), .C(_5181_), .Y(_5184_) );
	AOI22X1 AOI22X1_771 ( .A(_4938_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_5088_), .Y(_5185_) );
	AOI22X1 AOI22X1_772 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_4887_), .C(_4860_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_5186_) );
	INVX1 INVX1_624 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_5187_) );
	NAND2X1 NAND2X1_1003 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_4977_), .Y(_5188_) );
	OAI21X1 OAI21X1_163 ( .A(_5187_), .B(_4949_), .C(_5188_), .Y(_5189_) );
	INVX1 INVX1_625 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_5190_) );
	NAND2X1 NAND2X1_1004 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_4903_), .Y(_5191_) );
	OAI21X1 OAI21X1_164 ( .A(_5190_), .B(_4906_), .C(_5191_), .Y(_5192_) );
	NOR2X1 NOR2X1_582 ( .A(_5189_), .B(_5192_), .Y(_5193_) );
	NAND3X1 NAND3X1_241 ( .A(_5185_), .B(_5186_), .C(_5193_), .Y(_5194_) );
	INVX1 INVX1_626 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_5195_) );
	NAND2X1 NAND2X1_1005 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_4885_), .Y(_5196_) );
	OAI21X1 OAI21X1_165 ( .A(_5195_), .B(_4915_), .C(_5196_), .Y(_5197_) );
	INVX1 INVX1_627 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_5198_) );
	INVX1 INVX1_628 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_5199_) );
	OAI22X1 OAI22X1_132 ( .A(_5198_), .B(_4921_), .C(_4919_), .D(_5199_), .Y(_5200_) );
	NOR2X1 NOR2X1_583 ( .A(_5200_), .B(_5197_), .Y(_5201_) );
	AOI22X1 AOI22X1_773 ( .A(_5005_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_4978_), .Y(_5202_) );
	AND2X2 AND2X2_107 ( .A(_4877_), .B(_4899_), .Y(_5203_) );
	AOI22X1 AOI22X1_774 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_5203_), .C(_5107_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_5204_) );
	NAND3X1 NAND3X1_242 ( .A(_5202_), .B(_5204_), .C(_5201_), .Y(_5205_) );
	NOR3X1 NOR3X1_420 ( .A(_5205_), .B(_5184_), .C(_5194_), .Y(_5206_) );
	INVX1 INVX1_629 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_5207_) );
	NOR3X1 NOR3X1_421 ( .A(_5207_), .B(_4872_), .C(_4871_), .Y(_5208_) );
	AND2X2 AND2X2_108 ( .A(_4893_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_5209_) );
	AND2X2 AND2X2_109 ( .A(_5013_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_5210_) );
	NOR3X1 NOR3X1_422 ( .A(_5210_), .B(_5209_), .C(_5208_), .Y(_5211_) );
	INVX1 INVX1_630 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_5212_) );
	INVX1 INVX1_631 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_5213_) );
	OAI22X1 OAI22X1_133 ( .A(_5213_), .B(_4948_), .C(_4898_), .D(_5212_), .Y(_5214_) );
	INVX1 INVX1_632 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_5215_) );
	INVX1 INVX1_633 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_5216_) );
	NAND2X1 NAND2X1_1006 ( .A(_4889_), .B(_4890_), .Y(_5217_) );
	OAI22X1 OAI22X1_134 ( .A(_5217_), .B(_5216_), .C(_5215_), .D(_4868_), .Y(_5218_) );
	NOR2X1 NOR2X1_584 ( .A(_5214_), .B(_5218_), .Y(_5219_) );
	INVX1 INVX1_634 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_5220_) );
	NOR3X1 NOR3X1_423 ( .A(_4849_), .B(_4866_), .C(_4857_), .Y(_5221_) );
	NAND2X1 NAND2X1_1007 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_5221_), .Y(_5222_) );
	OAI21X1 OAI21X1_166 ( .A(_4878_), .B(_5220_), .C(_5222_), .Y(_5223_) );
	INVX1 INVX1_635 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_5224_) );
	INVX1 INVX1_636 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_5225_) );
	OAI22X1 OAI22X1_135 ( .A(_4965_), .B(_5225_), .C(_5224_), .D(_4966_), .Y(_5226_) );
	NOR2X1 NOR2X1_585 ( .A(_5223_), .B(_5226_), .Y(_5227_) );
	NAND3X1 NAND3X1_243 ( .A(_5211_), .B(_5227_), .C(_5219_), .Y(_5228_) );
	AOI22X1 AOI22X1_775 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_4970_), .C(_4971_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_5229_) );
	AOI22X1 AOI22X1_776 ( .A(_4973_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_4974_), .Y(_5230_) );
	NAND2X1 NAND2X1_1008 ( .A(_5229_), .B(_5230_), .Y(_5231_) );
	AOI22X1 AOI22X1_777 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_4981_), .C(_4980_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_5232_) );
	AOI22X1 AOI22X1_778 ( .A(_4924_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_4931_), .Y(_5233_) );
	NAND2X1 NAND2X1_1009 ( .A(_5232_), .B(_5233_), .Y(_5234_) );
	NOR2X1 NOR2X1_586 ( .A(_5231_), .B(_5234_), .Y(_5235_) );
	AOI22X1 AOI22X1_779 ( .A(_4985_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_4986_), .Y(_5236_) );
	AOI22X1 AOI22X1_780 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_5012_), .C(_4988_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_5237_) );
	NAND2X1 NAND2X1_1010 ( .A(_5237_), .B(_5236_), .Y(_5238_) );
	AOI22X1 AOI22X1_781 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_4992_), .C(_4993_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_5239_) );
	AOI22X1 AOI22X1_782 ( .A(_4995_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_4996_), .Y(_5240_) );
	NAND2X1 NAND2X1_1011 ( .A(_5240_), .B(_5239_), .Y(_5241_) );
	NOR2X1 NOR2X1_587 ( .A(_5238_), .B(_5241_), .Y(_5242_) );
	NAND2X1 NAND2X1_1012 ( .A(_5242_), .B(_5235_), .Y(_5243_) );
	AOI22X1 AOI22X1_783 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_5002_), .C(_5001_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_5244_) );
	AOI22X1 AOI22X1_784 ( .A(_4926_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_5004_), .Y(_5245_) );
	NAND2X1 NAND2X1_1013 ( .A(_5244_), .B(_5245_), .Y(_5246_) );
	AOI22X1 AOI22X1_785 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_5010_), .C(_5008_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_5247_) );
	AOI22X1 AOI22X1_786 ( .A(_4940_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_4958_), .Y(_5248_) );
	NAND2X1 NAND2X1_1014 ( .A(_5248_), .B(_5247_), .Y(_5249_) );
	NOR2X1 NOR2X1_588 ( .A(_5249_), .B(_5246_), .Y(_5250_) );
	AOI22X1 AOI22X1_787 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_5017_), .C(_5018_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_5251_) );
	NAND2X1 NAND2X1_1015 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_5020_), .Y(_5252_) );
	NAND2X1 NAND2X1_1016 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_5022_), .Y(_5253_) );
	NAND3X1 NAND3X1_244 ( .A(_5252_), .B(_5253_), .C(_5251_), .Y(_5254_) );
	AOI22X1 AOI22X1_788 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_5026_), .C(_5025_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_5255_) );
	AOI22X1 AOI22X1_789 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_5029_), .C(_5028_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_5256_) );
	NAND2X1 NAND2X1_1017 ( .A(_5255_), .B(_5256_), .Y(_5257_) );
	NOR2X1 NOR2X1_589 ( .A(_5257_), .B(_5254_), .Y(_5258_) );
	NAND2X1 NAND2X1_1018 ( .A(_5250_), .B(_5258_), .Y(_5259_) );
	NOR3X1 NOR3X1_424 ( .A(_5243_), .B(_5228_), .C(_5259_), .Y(_5260_) );
	AOI22X1 AOI22X1_790 ( .A(_5066_), .B(wData[42]), .C(wData[38]), .D(_5068_), .Y(_5261_) );
	AOI22X1 AOI22X1_791 ( .A(_5063_), .B(wData[46]), .C(_5070_), .D(wData[2]), .Y(_5262_) );
	NAND2X1 NAND2X1_1019 ( .A(_5261_), .B(_5262_), .Y(_5263_) );
	AOI21X1 AOI21X1_117 ( .A(wData[34]), .B(_5056_), .C(_5263_), .Y(_5264_) );
	INVX1 INVX1_637 ( .A(wData[50]), .Y(_5265_) );
	AOI22X1 AOI22X1_792 ( .A(_5076_), .B(wData[10]), .C(wData[14]), .D(_5077_), .Y(_5266_) );
	OAI21X1 OAI21X1_167 ( .A(_5265_), .B(_5075_), .C(_5266_), .Y(_5267_) );
	AOI22X1 AOI22X1_793 ( .A(_5039_), .B(wData[22]), .C(wData[18]), .D(_5042_), .Y(_5268_) );
	NAND2X1 NAND2X1_1020 ( .A(wData[26]), .B(_5046_), .Y(_5269_) );
	AOI22X1 AOI22X1_794 ( .A(_5052_), .B(wData[30]), .C(wData[6]), .D(_5050_), .Y(_5270_) );
	NAND3X1 NAND3X1_245 ( .A(_5269_), .B(_5270_), .C(_5268_), .Y(_5271_) );
	NOR2X1 NOR2X1_590 ( .A(_5267_), .B(_5271_), .Y(_5272_) );
	NAND2X1 NAND2X1_1021 ( .A(wData[58]), .B(_5059_), .Y(_5273_) );
	NAND2X1 NAND2X1_1022 ( .A(wData[54]), .B(_5060_), .Y(_5274_) );
	NAND2X1 NAND2X1_1023 ( .A(_5273_), .B(_5274_), .Y(_5275_) );
	AOI21X1 AOI21X1_118 ( .A(wData[62]), .B(_5062_), .C(_5275_), .Y(_5276_) );
	NAND3X1 NAND3X1_246 ( .A(_5264_), .B(_5276_), .C(_5272_), .Y(_5277_) );
	NOR2X1 NOR2X1_591 ( .A(_4844_), .B(_5277_), .Y(_5278_) );
	AOI21X1 AOI21X1_119 ( .A(_5206_), .B(_5260_), .C(_5278_), .Y(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_2_) );
	AOI21X1 AOI21X1_120 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_5088_), .C(_4845_), .Y(_5279_) );
	AOI22X1 AOI22X1_795 ( .A(_4860_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_5180_), .Y(_5280_) );
	AOI22X1 AOI22X1_796 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_5182_), .C(_4938_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_5281_) );
	NAND3X1 NAND3X1_247 ( .A(_5281_), .B(_5279_), .C(_5280_), .Y(_5282_) );
	AOI22X1 AOI22X1_797 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_4887_), .C(_4885_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_5283_) );
	AOI22X1 AOI22X1_798 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_4958_), .C(_5083_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_5284_) );
	INVX1 INVX1_638 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_5285_) );
	INVX1 INVX1_639 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_5286_) );
	OAI22X1 OAI22X1_136 ( .A(_5285_), .B(_4900_), .C(_4949_), .D(_5286_), .Y(_5287_) );
	INVX1 INVX1_640 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_5288_) );
	NAND2X1 NAND2X1_1024 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_5001_), .Y(_5289_) );
	OAI21X1 OAI21X1_168 ( .A(_5288_), .B(_4906_), .C(_5289_), .Y(_5290_) );
	NOR2X1 NOR2X1_592 ( .A(_5287_), .B(_5290_), .Y(_5291_) );
	NAND3X1 NAND3X1_248 ( .A(_5283_), .B(_5284_), .C(_5291_), .Y(_5292_) );
	AND2X2 AND2X2_110 ( .A(_4914_), .B(_4848_), .Y(_5293_) );
	AOI22X1 AOI22X1_799 ( .A(_4853_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_5293_), .Y(_5294_) );
	AND2X2 AND2X2_111 ( .A(_4912_), .B(_4877_), .Y(_5295_) );
	AND2X2 AND2X2_112 ( .A(_4920_), .B(_4877_), .Y(_5296_) );
	AOI22X1 AOI22X1_800 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_5296_), .C(_5295_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_5297_) );
	NAND2X1 NAND2X1_1025 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_5005_), .Y(_5298_) );
	NAND2X1 NAND2X1_1026 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_4978_), .Y(_5299_) );
	NAND2X1 NAND2X1_1027 ( .A(_5298_), .B(_5299_), .Y(_5300_) );
	INVX1 INVX1_641 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_5301_) );
	NAND2X1 NAND2X1_1028 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_4977_), .Y(_5302_) );
	OAI21X1 OAI21X1_169 ( .A(_5301_), .B(_4930_), .C(_5302_), .Y(_5303_) );
	NOR2X1 NOR2X1_593 ( .A(_5300_), .B(_5303_), .Y(_5304_) );
	NAND3X1 NAND3X1_249 ( .A(_5294_), .B(_5297_), .C(_5304_), .Y(_5305_) );
	NOR3X1 NOR3X1_425 ( .A(_5292_), .B(_5282_), .C(_5305_), .Y(_5306_) );
	INVX1 INVX1_642 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_5307_) );
	NAND2X1 NAND2X1_1029 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_4893_), .Y(_5308_) );
	OAI21X1 OAI21X1_170 ( .A(_4898_), .B(_5307_), .C(_5308_), .Y(_5309_) );
	AOI21X1 AOI21X1_121 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_4873_), .C(_5309_), .Y(_5310_) );
	INVX1 INVX1_643 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_5311_) );
	INVX1 INVX1_644 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_5312_) );
	OAI22X1 OAI22X1_137 ( .A(_5217_), .B(_5312_), .C(_5311_), .D(_4868_), .Y(_5313_) );
	INVX1 INVX1_645 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_5314_) );
	NAND2X1 NAND2X1_1030 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_5013_), .Y(_5315_) );
	OAI21X1 OAI21X1_171 ( .A(_4878_), .B(_5314_), .C(_5315_), .Y(_5316_) );
	NOR2X1 NOR2X1_594 ( .A(_5316_), .B(_5313_), .Y(_5317_) );
	INVX1 INVX1_646 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_5318_) );
	INVX1 INVX1_647 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_5319_) );
	OAI22X1 OAI22X1_138 ( .A(_4965_), .B(_5319_), .C(_5318_), .D(_4966_), .Y(_5320_) );
	INVX1 INVX1_648 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_5321_) );
	NAND2X1 NAND2X1_1031 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_5012_), .Y(_5322_) );
	OAI21X1 OAI21X1_172 ( .A(_5321_), .B(_4948_), .C(_5322_), .Y(_5323_) );
	NOR2X1 NOR2X1_595 ( .A(_5323_), .B(_5320_), .Y(_5324_) );
	NAND3X1 NAND3X1_250 ( .A(_5310_), .B(_5324_), .C(_5317_), .Y(_5325_) );
	AOI22X1 AOI22X1_801 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_4970_), .C(_4971_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_5326_) );
	AOI22X1 AOI22X1_802 ( .A(_4973_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_4974_), .Y(_5327_) );
	NAND2X1 NAND2X1_1032 ( .A(_5326_), .B(_5327_), .Y(_5328_) );
	AOI22X1 AOI22X1_803 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_4981_), .C(_4980_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_5329_) );
	AOI22X1 AOI22X1_804 ( .A(_4924_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_4931_), .Y(_5330_) );
	NAND2X1 NAND2X1_1033 ( .A(_5329_), .B(_5330_), .Y(_5331_) );
	NOR2X1 NOR2X1_596 ( .A(_5328_), .B(_5331_), .Y(_5332_) );
	AOI22X1 AOI22X1_805 ( .A(_4985_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_4986_), .Y(_5333_) );
	AOI22X1 AOI22X1_806 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_5221_), .C(_4988_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_5334_) );
	NAND2X1 NAND2X1_1034 ( .A(_5334_), .B(_5333_), .Y(_5335_) );
	AOI22X1 AOI22X1_807 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_4992_), .C(_4993_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_5336_) );
	AOI22X1 AOI22X1_808 ( .A(_4995_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_4996_), .Y(_5337_) );
	NAND2X1 NAND2X1_1035 ( .A(_5337_), .B(_5336_), .Y(_5338_) );
	NOR2X1 NOR2X1_597 ( .A(_5335_), .B(_5338_), .Y(_5339_) );
	NAND2X1 NAND2X1_1036 ( .A(_5339_), .B(_5332_), .Y(_5340_) );
	AOI22X1 AOI22X1_809 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_5002_), .C(_4903_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_5341_) );
	AOI22X1 AOI22X1_810 ( .A(_4926_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_5004_), .Y(_5342_) );
	NAND2X1 NAND2X1_1037 ( .A(_5341_), .B(_5342_), .Y(_5343_) );
	AOI22X1 AOI22X1_811 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_5010_), .C(_5008_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_5344_) );
	AOI22X1 AOI22X1_812 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_4940_), .C(_4989_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_5345_) );
	NAND2X1 NAND2X1_1038 ( .A(_5345_), .B(_5344_), .Y(_5346_) );
	NOR2X1 NOR2X1_598 ( .A(_5346_), .B(_5343_), .Y(_5347_) );
	AOI22X1 AOI22X1_813 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_5017_), .C(_5018_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_5348_) );
	NAND2X1 NAND2X1_1039 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_5020_), .Y(_5349_) );
	NAND2X1 NAND2X1_1040 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_5022_), .Y(_5350_) );
	NAND3X1 NAND3X1_251 ( .A(_5349_), .B(_5350_), .C(_5348_), .Y(_5351_) );
	AOI22X1 AOI22X1_814 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_5026_), .C(_5025_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_5352_) );
	AOI22X1 AOI22X1_815 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_5029_), .C(_5028_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_5353_) );
	NAND2X1 NAND2X1_1041 ( .A(_5352_), .B(_5353_), .Y(_5354_) );
	NOR2X1 NOR2X1_599 ( .A(_5354_), .B(_5351_), .Y(_5355_) );
	NAND2X1 NAND2X1_1042 ( .A(_5347_), .B(_5355_), .Y(_5356_) );
	NOR3X1 NOR3X1_426 ( .A(_5340_), .B(_5325_), .C(_5356_), .Y(_5357_) );
	NAND2X1 NAND2X1_1043 ( .A(wData[59]), .B(_5059_), .Y(_5358_) );
	OAI21X1 OAI21X1_173 ( .A(_4843_), .B(wBusy_bF_buf3), .C(_5358_), .Y(_5359_) );
	NAND2X1 NAND2X1_1044 ( .A(wData[7]), .B(_5050_), .Y(_5360_) );
	NAND2X1 NAND2X1_1045 ( .A(wData[55]), .B(_5060_), .Y(_5361_) );
	AOI22X1 AOI22X1_816 ( .A(wData[63]), .B(_5062_), .C(_5052_), .D(wData[31]), .Y(_5362_) );
	NAND3X1 NAND3X1_252 ( .A(_5360_), .B(_5361_), .C(_5362_), .Y(_5363_) );
	OR2X2 OR2X2_57 ( .A(_5363_), .B(_5359_), .Y(_5364_) );
	INVX1 INVX1_649 ( .A(wData[51]), .Y(_5365_) );
	NAND2X1 NAND2X1_1046 ( .A(wData[47]), .B(_5063_), .Y(_5366_) );
	OAI21X1 OAI21X1_174 ( .A(_5365_), .B(_5075_), .C(_5366_), .Y(_5367_) );
	AOI21X1 AOI21X1_122 ( .A(wData[3]), .B(_5070_), .C(_5367_), .Y(_5368_) );
	AOI22X1 AOI22X1_817 ( .A(_5076_), .B(wData[11]), .C(wData[15]), .D(_5077_), .Y(_5369_) );
	AOI22X1 AOI22X1_818 ( .A(_5039_), .B(wData[23]), .C(wData[27]), .D(_5046_), .Y(_5370_) );
	AND2X2 AND2X2_113 ( .A(_5369_), .B(_5370_), .Y(_5371_) );
	NAND2X1 NAND2X1_1047 ( .A(wData[39]), .B(_5068_), .Y(_5372_) );
	NAND2X1 NAND2X1_1048 ( .A(wData[43]), .B(_5066_), .Y(_5373_) );
	NAND2X1 NAND2X1_1049 ( .A(_5372_), .B(_5373_), .Y(_5374_) );
	NAND2X1 NAND2X1_1050 ( .A(wData[19]), .B(_5042_), .Y(_5375_) );
	NAND2X1 NAND2X1_1051 ( .A(wData[35]), .B(_5056_), .Y(_5376_) );
	NAND2X1 NAND2X1_1052 ( .A(_5375_), .B(_5376_), .Y(_5377_) );
	NOR2X1 NOR2X1_600 ( .A(_5374_), .B(_5377_), .Y(_5378_) );
	NAND3X1 NAND3X1_253 ( .A(_5371_), .B(_5368_), .C(_5378_), .Y(_5379_) );
	NOR2X1 NOR2X1_601 ( .A(_5364_), .B(_5379_), .Y(_5380_) );
	AOI21X1 AOI21X1_123 ( .A(_5306_), .B(_5357_), .C(_5380_), .Y(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_3_) );
	INVX1 INVX1_650 ( .A(wSelec[110]), .Y(_5381_) );
	NOR2X1 NOR2X1_602 ( .A(wBusy_bF_buf2), .B(_5381_), .Y(_5382_) );
	INVX1 INVX1_651 ( .A(_5382_), .Y(_5383_) );
	INVX1 INVX1_652 ( .A(wSelec[120]), .Y(_5384_) );
	NAND2X1 NAND2X1_1053 ( .A(wSelec[119]), .B(_5384_), .Y(_5385_) );
	INVX2 INVX2_17 ( .A(_5385_), .Y(_5386_) );
	OR2X2 OR2X2_58 ( .A(wSelec[116]), .B(wSelec[115]), .Y(_5387_) );
	INVX1 INVX1_653 ( .A(wSelec[118]), .Y(_5388_) );
	NAND2X1 NAND2X1_1054 ( .A(wSelec[117]), .B(_5388_), .Y(_5389_) );
	NOR2X1 NOR2X1_603 ( .A(_5387_), .B(_5389_), .Y(_5390_) );
	AND2X2 AND2X2_114 ( .A(_5390_), .B(_5386_), .Y(_5391_) );
	AOI21X1 AOI21X1_124 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_5391_), .C(_5383_), .Y(_5392_) );
	INVX1 INVX1_654 ( .A(wSelec[116]), .Y(_5393_) );
	NAND2X1 NAND2X1_1055 ( .A(wSelec[115]), .B(_5393_), .Y(_5394_) );
	OR2X2 OR2X2_59 ( .A(wSelec[117]), .B(wSelec[118]), .Y(_5395_) );
	NOR2X1 NOR2X1_604 ( .A(_5395_), .B(_5394_), .Y(_5396_) );
	NAND2X1 NAND2X1_1056 ( .A(_5386_), .B(_5396_), .Y(_5397_) );
	INVX1 INVX1_655 ( .A(_5397_), .Y(_5398_) );
	INVX1 INVX1_656 ( .A(wSelec[115]), .Y(_5399_) );
	NAND2X1 NAND2X1_1057 ( .A(wSelec[116]), .B(_5399_), .Y(_5400_) );
	INVX1 INVX1_657 ( .A(wSelec[117]), .Y(_5401_) );
	NAND2X1 NAND2X1_1058 ( .A(wSelec[118]), .B(_5401_), .Y(_5402_) );
	NOR2X1 NOR2X1_605 ( .A(_5400_), .B(_5402_), .Y(_5403_) );
	NAND2X1 NAND2X1_1059 ( .A(wSelec[119]), .B(wSelec[120]), .Y(_5404_) );
	INVX1 INVX1_658 ( .A(_5404_), .Y(_5405_) );
	NAND2X1 NAND2X1_1060 ( .A(_5405_), .B(_5403_), .Y(_5406_) );
	INVX1 INVX1_659 ( .A(_5406_), .Y(_5407_) );
	AOI22X1 AOI22X1_819 ( .A(_5398_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_5407_), .Y(_5408_) );
	OR2X2 OR2X2_60 ( .A(_5394_), .B(_5395_), .Y(_5409_) );
	OR2X2 OR2X2_61 ( .A(wSelec[119]), .B(wSelec[120]), .Y(_5410_) );
	NOR2X1 NOR2X1_606 ( .A(_5410_), .B(_5409_), .Y(_5411_) );
	NOR2X1 NOR2X1_607 ( .A(_5389_), .B(_5394_), .Y(_5412_) );
	INVX1 INVX1_660 ( .A(wSelec[119]), .Y(_5413_) );
	NAND2X1 NAND2X1_1061 ( .A(wSelec[120]), .B(_5413_), .Y(_5414_) );
	INVX2 INVX2_18 ( .A(_5414_), .Y(_5415_) );
	NAND2X1 NAND2X1_1062 ( .A(_5415_), .B(_5412_), .Y(_5416_) );
	INVX1 INVX1_661 ( .A(_5416_), .Y(_5417_) );
	AOI22X1 AOI22X1_820 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_5411_), .C(_5417_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_5418_) );
	NAND3X1 NAND3X1_254 ( .A(_5392_), .B(_5418_), .C(_5408_), .Y(_5419_) );
	NOR2X1 NOR2X1_608 ( .A(wSelec[116]), .B(wSelec[115]), .Y(_5420_) );
	NOR2X1 NOR2X1_609 ( .A(wSelec[117]), .B(wSelec[118]), .Y(_5421_) );
	NAND2X1 NAND2X1_1063 ( .A(_5420_), .B(_5421_), .Y(_5422_) );
	NOR2X1 NOR2X1_610 ( .A(_5385_), .B(_5422_), .Y(_5423_) );
	NAND2X1 NAND2X1_1064 ( .A(wSelec[116]), .B(wSelec[115]), .Y(_5424_) );
	NOR3X1 NOR3X1_427 ( .A(_5395_), .B(_5424_), .C(_5385_), .Y(_5425_) );
	AOI22X1 AOI22X1_821 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_5425_), .C(_5423_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_5426_) );
	INVX1 INVX1_662 ( .A(_5410_), .Y(_5427_) );
	NOR2X1 NOR2X1_611 ( .A(_5395_), .B(_5400_), .Y(_5428_) );
	AND2X2 AND2X2_115 ( .A(_5428_), .B(_5427_), .Y(_5429_) );
	NAND2X1 NAND2X1_1065 ( .A(wSelec[117]), .B(wSelec[118]), .Y(_5430_) );
	NOR3X1 NOR3X1_428 ( .A(_5404_), .B(_5424_), .C(_5430_), .Y(_5431_) );
	AOI22X1 AOI22X1_822 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_5431_), .C(_5429_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_5432_) );
	INVX1 INVX1_663 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_5433_) );
	INVX1 INVX1_664 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_5434_) );
	NOR2X1 NOR2X1_612 ( .A(_5394_), .B(_5402_), .Y(_5435_) );
	NAND2X1 NAND2X1_1066 ( .A(_5405_), .B(_5435_), .Y(_5436_) );
	NOR2X1 NOR2X1_613 ( .A(_5424_), .B(_5430_), .Y(_5437_) );
	NAND2X1 NAND2X1_1067 ( .A(_5437_), .B(_5415_), .Y(_5438_) );
	OAI22X1 OAI22X1_139 ( .A(_5433_), .B(_5438_), .C(_5436_), .D(_5434_), .Y(_5439_) );
	INVX1 INVX1_665 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_5440_) );
	NOR3X1 NOR3X1_429 ( .A(_5385_), .B(_5400_), .C(_5402_), .Y(_5441_) );
	NAND2X1 NAND2X1_1068 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_5441_), .Y(_5442_) );
	NOR2X1 NOR2X1_614 ( .A(_5424_), .B(_5389_), .Y(_5443_) );
	NAND2X1 NAND2X1_1069 ( .A(_5415_), .B(_5443_), .Y(_5444_) );
	OAI21X1 OAI21X1_175 ( .A(_5440_), .B(_5444_), .C(_5442_), .Y(_5445_) );
	NOR2X1 NOR2X1_615 ( .A(_5439_), .B(_5445_), .Y(_5446_) );
	NAND3X1 NAND3X1_255 ( .A(_5426_), .B(_5432_), .C(_5446_), .Y(_5447_) );
	INVX1 INVX1_666 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_5448_) );
	INVX1 INVX1_667 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_5449_) );
	NOR2X1 NOR2X1_616 ( .A(_5389_), .B(_5400_), .Y(_5450_) );
	NAND2X1 NAND2X1_1070 ( .A(_5386_), .B(_5450_), .Y(_5451_) );
	NOR2X1 NOR2X1_617 ( .A(_5387_), .B(_5402_), .Y(_5452_) );
	NAND2X1 NAND2X1_1071 ( .A(_5386_), .B(_5452_), .Y(_5453_) );
	OAI22X1 OAI22X1_140 ( .A(_5453_), .B(_5448_), .C(_5449_), .D(_5451_), .Y(_5454_) );
	INVX1 INVX1_668 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_5455_) );
	INVX1 INVX1_669 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_5456_) );
	NAND2X1 NAND2X1_1072 ( .A(_5415_), .B(_5450_), .Y(_5457_) );
	NOR2X1 NOR2X1_618 ( .A(_5424_), .B(_5395_), .Y(_5458_) );
	NAND2X1 NAND2X1_1073 ( .A(_5415_), .B(_5458_), .Y(_5459_) );
	OAI22X1 OAI22X1_141 ( .A(_5455_), .B(_5459_), .C(_5457_), .D(_5456_), .Y(_5460_) );
	NOR2X1 NOR2X1_619 ( .A(_5460_), .B(_5454_), .Y(_5461_) );
	NOR3X1 NOR3X1_430 ( .A(_5394_), .B(_5430_), .C(_5414_), .Y(_5462_) );
	NAND2X1 NAND2X1_1074 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_5462_), .Y(_5463_) );
	NOR3X1 NOR3X1_431 ( .A(_5402_), .B(_5424_), .C(_5414_), .Y(_5464_) );
	NAND2X1 NAND2X1_1075 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_5464_), .Y(_5465_) );
	NAND2X1 NAND2X1_1076 ( .A(_5463_), .B(_5465_), .Y(_5466_) );
	INVX1 INVX1_670 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_5467_) );
	NAND2X1 NAND2X1_1077 ( .A(_5405_), .B(_5390_), .Y(_5468_) );
	NOR3X1 NOR3X1_432 ( .A(_5400_), .B(_5402_), .C(_5414_), .Y(_5469_) );
	NAND2X1 NAND2X1_1078 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_5469_), .Y(_5470_) );
	OAI21X1 OAI21X1_176 ( .A(_5467_), .B(_5468_), .C(_5470_), .Y(_5471_) );
	NOR2X1 NOR2X1_620 ( .A(_5466_), .B(_5471_), .Y(_5472_) );
	NAND2X1 NAND2X1_1079 ( .A(_5461_), .B(_5472_), .Y(_5473_) );
	NOR3X1 NOR3X1_433 ( .A(_5419_), .B(_5473_), .C(_5447_), .Y(_5474_) );
	NAND2X1 NAND2X1_1080 ( .A(_5386_), .B(_5443_), .Y(_5475_) );
	INVX1 INVX1_671 ( .A(_5475_), .Y(_5476_) );
	INVX1 INVX1_672 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_5477_) );
	NOR3X1 NOR3X1_434 ( .A(_5387_), .B(_5410_), .C(_5389_), .Y(_5478_) );
	NAND2X1 NAND2X1_1081 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_5478_), .Y(_5479_) );
	NAND2X1 NAND2X1_1082 ( .A(_5427_), .B(_5450_), .Y(_5480_) );
	OAI21X1 OAI21X1_177 ( .A(_5480_), .B(_5477_), .C(_5479_), .Y(_5481_) );
	AOI21X1 AOI21X1_125 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_5476_), .C(_5481_), .Y(_5482_) );
	INVX1 INVX1_673 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_5483_) );
	INVX1 INVX1_674 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_5484_) );
	NOR2X1 NOR2X1_621 ( .A(_5430_), .B(_5387_), .Y(_5485_) );
	NAND2X1 NAND2X1_1083 ( .A(_5386_), .B(_5485_), .Y(_5486_) );
	NAND2X1 NAND2X1_1084 ( .A(_5427_), .B(_5412_), .Y(_5487_) );
	OAI22X1 OAI22X1_142 ( .A(_5484_), .B(_5486_), .C(_5487_), .D(_5483_), .Y(_5488_) );
	INVX1 INVX1_675 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_5489_) );
	INVX1 INVX1_676 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_5490_) );
	NAND2X1 NAND2X1_1085 ( .A(_5386_), .B(_5412_), .Y(_5491_) );
	NAND2X1 NAND2X1_1086 ( .A(_5427_), .B(_5458_), .Y(_5492_) );
	OAI22X1 OAI22X1_143 ( .A(_5489_), .B(_5492_), .C(_5491_), .D(_5490_), .Y(_5493_) );
	NOR2X1 NOR2X1_622 ( .A(_5488_), .B(_5493_), .Y(_5494_) );
	INVX1 INVX1_677 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_5495_) );
	NOR3X1 NOR3X1_435 ( .A(_5410_), .B(_5424_), .C(_5389_), .Y(_5496_) );
	NAND2X1 NAND2X1_1087 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_5496_), .Y(_5497_) );
	OR2X2 OR2X2_62 ( .A(_5422_), .B(_5404_), .Y(_5498_) );
	OAI21X1 OAI21X1_178 ( .A(_5495_), .B(_5498_), .C(_5497_), .Y(_5499_) );
	INVX1 INVX1_678 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_5500_) );
	INVX1 INVX1_679 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_5501_) );
	NOR2X1 NOR2X1_623 ( .A(_5430_), .B(_5400_), .Y(_5502_) );
	NAND2X1 NAND2X1_1088 ( .A(_5386_), .B(_5502_), .Y(_5503_) );
	NAND2X1 NAND2X1_1089 ( .A(_5405_), .B(_5396_), .Y(_5504_) );
	OAI22X1 OAI22X1_144 ( .A(_5503_), .B(_5501_), .C(_5500_), .D(_5504_), .Y(_5505_) );
	NOR2X1 NOR2X1_624 ( .A(_5499_), .B(_5505_), .Y(_5506_) );
	NAND3X1 NAND3X1_256 ( .A(_5482_), .B(_5506_), .C(_5494_), .Y(_5507_) );
	NOR3X1 NOR3X1_436 ( .A(_5387_), .B(_5395_), .C(_5410_), .Y(_5508_) );
	NOR3X1 NOR3X1_437 ( .A(_5404_), .B(_5430_), .C(_5394_), .Y(_5509_) );
	AOI22X1 AOI22X1_823 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_5508_), .C(_5509_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_5510_) );
	NOR3X1 NOR3X1_438 ( .A(_5404_), .B(_5430_), .C(_5400_), .Y(_5511_) );
	NOR3X1 NOR3X1_439 ( .A(_5404_), .B(_5424_), .C(_5402_), .Y(_5512_) );
	AOI22X1 AOI22X1_824 ( .A(_5511_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_5512_), .Y(_5513_) );
	NAND2X1 NAND2X1_1090 ( .A(_5510_), .B(_5513_), .Y(_5514_) );
	NOR3X1 NOR3X1_440 ( .A(_5402_), .B(_5387_), .C(_5414_), .Y(_5515_) );
	NOR3X1 NOR3X1_441 ( .A(_5394_), .B(_5402_), .C(_5414_), .Y(_5516_) );
	AOI22X1 AOI22X1_825 ( .A(_5515_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_5516_), .Y(_5517_) );
	NOR3X1 NOR3X1_442 ( .A(_5385_), .B(_5430_), .C(_5394_), .Y(_5518_) );
	NOR3X1 NOR3X1_443 ( .A(_5424_), .B(_5430_), .C(_5385_), .Y(_5519_) );
	AOI22X1 AOI22X1_826 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_5519_), .C(_5518_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_5520_) );
	NAND2X1 NAND2X1_1091 ( .A(_5520_), .B(_5517_), .Y(_5521_) );
	NOR2X1 NOR2X1_625 ( .A(_5514_), .B(_5521_), .Y(_5522_) );
	NOR3X1 NOR3X1_444 ( .A(_5410_), .B(_5430_), .C(_5394_), .Y(_5523_) );
	NOR3X1 NOR3X1_445 ( .A(_5410_), .B(_5430_), .C(_5400_), .Y(_5524_) );
	AOI22X1 AOI22X1_827 ( .A(_5523_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_5524_), .Y(_5525_) );
	NOR3X1 NOR3X1_446 ( .A(_5410_), .B(_5424_), .C(_5402_), .Y(_5526_) );
	NOR3X1 NOR3X1_447 ( .A(_5385_), .B(_5395_), .C(_5400_), .Y(_5527_) );
	AOI22X1 AOI22X1_828 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_5526_), .C(_5527_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_5528_) );
	NAND2X1 NAND2X1_1092 ( .A(_5525_), .B(_5528_), .Y(_5529_) );
	NOR3X1 NOR3X1_448 ( .A(_5424_), .B(_5430_), .C(_5410_), .Y(_5530_) );
	NOR3X1 NOR3X1_449 ( .A(_5400_), .B(_5395_), .C(_5414_), .Y(_5531_) );
	AOI22X1 AOI22X1_829 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_5530_), .C(_5531_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_5532_) );
	NOR3X1 NOR3X1_450 ( .A(_5387_), .B(_5395_), .C(_5414_), .Y(_5533_) );
	NOR3X1 NOR3X1_451 ( .A(_5387_), .B(_5430_), .C(_5414_), .Y(_5534_) );
	AOI22X1 AOI22X1_830 ( .A(_5533_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_5534_), .Y(_5535_) );
	NAND2X1 NAND2X1_1093 ( .A(_5535_), .B(_5532_), .Y(_5536_) );
	NOR2X1 NOR2X1_626 ( .A(_5529_), .B(_5536_), .Y(_5537_) );
	NAND2X1 NAND2X1_1094 ( .A(_5537_), .B(_5522_), .Y(_5538_) );
	NOR3X1 NOR3X1_452 ( .A(_5385_), .B(_5424_), .C(_5402_), .Y(_5539_) );
	NOR3X1 NOR3X1_453 ( .A(_5395_), .B(_5404_), .C(_5400_), .Y(_5540_) );
	AOI22X1 AOI22X1_831 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_5540_), .C(_5539_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_5541_) );
	NOR3X1 NOR3X1_454 ( .A(_5389_), .B(_5387_), .C(_5414_), .Y(_5542_) );
	NOR3X1 NOR3X1_455 ( .A(_5400_), .B(_5430_), .C(_5414_), .Y(_5543_) );
	AOI22X1 AOI22X1_832 ( .A(_5542_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_5543_), .Y(_5544_) );
	NAND2X1 NAND2X1_1095 ( .A(_5541_), .B(_5544_), .Y(_5545_) );
	NOR3X1 NOR3X1_456 ( .A(_5385_), .B(_5394_), .C(_5402_), .Y(_5546_) );
	NAND2X1 NAND2X1_1096 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_5546_), .Y(_5547_) );
	NOR3X1 NOR3X1_457 ( .A(_5404_), .B(_5424_), .C(_5389_), .Y(_5548_) );
	NAND2X1 NAND2X1_1097 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_5548_), .Y(_5549_) );
	NOR3X1 NOR3X1_458 ( .A(_5387_), .B(_5430_), .C(_5410_), .Y(_5550_) );
	NOR3X1 NOR3X1_459 ( .A(_5387_), .B(_5404_), .C(_5402_), .Y(_5551_) );
	AOI22X1 AOI22X1_833 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_5550_), .C(_5551_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_5552_) );
	NAND3X1 NAND3X1_257 ( .A(_5547_), .B(_5549_), .C(_5552_), .Y(_5553_) );
	NOR2X1 NOR2X1_627 ( .A(_5553_), .B(_5545_), .Y(_5554_) );
	NOR3X1 NOR3X1_460 ( .A(_5387_), .B(_5410_), .C(_5402_), .Y(_5555_) );
	NOR3X1 NOR3X1_461 ( .A(_5389_), .B(_5404_), .C(_5394_), .Y(_5556_) );
	AOI22X1 AOI22X1_834 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_5555_), .C(_5556_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_5557_) );
	NOR3X1 NOR3X1_462 ( .A(_5389_), .B(_5404_), .C(_5400_), .Y(_5558_) );
	NAND2X1 NAND2X1_1098 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_5558_), .Y(_5559_) );
	NOR3X1 NOR3X1_463 ( .A(_5394_), .B(_5395_), .C(_5414_), .Y(_5560_) );
	NAND2X1 NAND2X1_1099 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_5560_), .Y(_5561_) );
	NAND3X1 NAND3X1_258 ( .A(_5559_), .B(_5561_), .C(_5557_), .Y(_5562_) );
	NOR3X1 NOR3X1_464 ( .A(_5394_), .B(_5410_), .C(_5402_), .Y(_5563_) );
	NOR3X1 NOR3X1_465 ( .A(_5404_), .B(_5430_), .C(_5387_), .Y(_5564_) );
	AOI22X1 AOI22X1_835 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_5564_), .C(_5563_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_5565_) );
	NOR3X1 NOR3X1_466 ( .A(_5400_), .B(_5410_), .C(_5402_), .Y(_5566_) );
	NOR3X1 NOR3X1_467 ( .A(_5404_), .B(_5424_), .C(_5395_), .Y(_5567_) );
	AOI22X1 AOI22X1_836 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_5567_), .C(_5566_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_5568_) );
	NAND2X1 NAND2X1_1100 ( .A(_5565_), .B(_5568_), .Y(_5569_) );
	NOR2X1 NOR2X1_628 ( .A(_5569_), .B(_5562_), .Y(_5570_) );
	NAND2X1 NAND2X1_1101 ( .A(_5554_), .B(_5570_), .Y(_5571_) );
	NOR3X1 NOR3X1_468 ( .A(_5538_), .B(_5507_), .C(_5571_), .Y(_5572_) );
	INVX1 INVX1_680 ( .A(wSelec[112]), .Y(_5573_) );
	NAND2X1 NAND2X1_1102 ( .A(wSelec[111]), .B(_5573_), .Y(_5574_) );
	INVX1 INVX1_681 ( .A(wSelec[114]), .Y(_5575_) );
	NAND2X1 NAND2X1_1103 ( .A(wSelec[113]), .B(_5575_), .Y(_5576_) );
	NOR2X1 NOR2X1_629 ( .A(_5574_), .B(_5576_), .Y(_5577_) );
	NOR2X1 NOR2X1_630 ( .A(wSelec[112]), .B(wSelec[111]), .Y(_5578_) );
	INVX1 INVX1_682 ( .A(_5578_), .Y(_5579_) );
	NOR2X1 NOR2X1_631 ( .A(_5576_), .B(_5579_), .Y(_5580_) );
	AOI22X1 AOI22X1_837 ( .A(wData[20]), .B(_5577_), .C(_5580_), .D(wData[16]), .Y(_5581_) );
	INVX1 INVX1_683 ( .A(wSelec[111]), .Y(_5582_) );
	NAND2X1 NAND2X1_1104 ( .A(wSelec[112]), .B(_5582_), .Y(_5583_) );
	NOR2X1 NOR2X1_632 ( .A(_5583_), .B(_5576_), .Y(_5584_) );
	NAND2X1 NAND2X1_1105 ( .A(wData[24]), .B(_5584_), .Y(_5585_) );
	INVX1 INVX1_684 ( .A(wSelec[113]), .Y(_5586_) );
	NAND2X1 NAND2X1_1106 ( .A(_5586_), .B(_5575_), .Y(_5587_) );
	NOR2X1 NOR2X1_633 ( .A(_5574_), .B(_5587_), .Y(_5588_) );
	NAND2X1 NAND2X1_1107 ( .A(wSelec[112]), .B(wSelec[111]), .Y(_5589_) );
	NOR2X1 NOR2X1_634 ( .A(_5589_), .B(_5576_), .Y(_5590_) );
	AOI22X1 AOI22X1_838 ( .A(_5590_), .B(wData[28]), .C(wData[4]), .D(_5588_), .Y(_5591_) );
	NAND3X1 NAND3X1_259 ( .A(_5585_), .B(_5591_), .C(_5581_), .Y(_5592_) );
	NAND2X1 NAND2X1_1108 ( .A(wSelec[114]), .B(_5586_), .Y(_5593_) );
	NOR2X1 NOR2X1_635 ( .A(_5593_), .B(_5579_), .Y(_5594_) );
	NAND2X1 NAND2X1_1109 ( .A(wData[32]), .B(_5594_), .Y(_5595_) );
	NAND2X1 NAND2X1_1110 ( .A(wSelec[113]), .B(wSelec[114]), .Y(_5596_) );
	NOR2X1 NOR2X1_636 ( .A(_5596_), .B(_5583_), .Y(_5597_) );
	NOR2X1 NOR2X1_637 ( .A(_5596_), .B(_5574_), .Y(_5598_) );
	AOI22X1 AOI22X1_839 ( .A(_5597_), .B(wData[56]), .C(wData[52]), .D(_5598_), .Y(_5599_) );
	NOR2X1 NOR2X1_638 ( .A(_5589_), .B(_5596_), .Y(_5600_) );
	NOR2X1 NOR2X1_639 ( .A(_5589_), .B(_5593_), .Y(_5601_) );
	AOI22X1 AOI22X1_840 ( .A(wData[60]), .B(_5600_), .C(_5601_), .D(wData[44]), .Y(_5602_) );
	NAND3X1 NAND3X1_260 ( .A(_5595_), .B(_5602_), .C(_5599_), .Y(_5603_) );
	NOR2X1 NOR2X1_640 ( .A(_5583_), .B(_5593_), .Y(_5604_) );
	NAND2X1 NAND2X1_1111 ( .A(wData[40]), .B(_5604_), .Y(_5605_) );
	NOR2X1 NOR2X1_641 ( .A(_5593_), .B(_5574_), .Y(_5606_) );
	NAND2X1 NAND2X1_1112 ( .A(wData[36]), .B(_5606_), .Y(_5607_) );
	NOR2X1 NOR2X1_642 ( .A(_5587_), .B(_5579_), .Y(_5608_) );
	NAND2X1 NAND2X1_1113 ( .A(wData[0]), .B(_5608_), .Y(_5609_) );
	NAND3X1 NAND3X1_261 ( .A(_5605_), .B(_5607_), .C(_5609_), .Y(_5610_) );
	INVX1 INVX1_685 ( .A(wData[48]), .Y(_5611_) );
	NOR2X1 NOR2X1_643 ( .A(_5586_), .B(_5575_), .Y(_5612_) );
	NAND2X1 NAND2X1_1114 ( .A(_5578_), .B(_5612_), .Y(_5613_) );
	NOR2X1 NOR2X1_644 ( .A(_5583_), .B(_5587_), .Y(_5614_) );
	NOR2X1 NOR2X1_645 ( .A(_5589_), .B(_5587_), .Y(_5615_) );
	AOI22X1 AOI22X1_841 ( .A(_5614_), .B(wData[8]), .C(wData[12]), .D(_5615_), .Y(_5616_) );
	OAI21X1 OAI21X1_179 ( .A(_5611_), .B(_5613_), .C(_5616_), .Y(_5617_) );
	OR2X2 OR2X2_63 ( .A(_5617_), .B(_5610_), .Y(_5618_) );
	NOR3X1 NOR3X1_469 ( .A(_5592_), .B(_5603_), .C(_5618_), .Y(_5619_) );
	AND2X2 AND2X2_116 ( .A(_5619_), .B(_5383_), .Y(_5620_) );
	AOI21X1 AOI21X1_126 ( .A(_5474_), .B(_5572_), .C(_5620_), .Y(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_0_) );
	INVX1 INVX1_686 ( .A(_5491_), .Y(_5621_) );
	AOI21X1 AOI21X1_127 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_5621_), .C(_5383_), .Y(_5622_) );
	AOI22X1 AOI22X1_842 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_5391_), .C(_5407_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_5623_) );
	AOI22X1 AOI22X1_843 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_5411_), .C(_5417_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_5624_) );
	NAND3X1 NAND3X1_262 ( .A(_5622_), .B(_5623_), .C(_5624_), .Y(_5625_) );
	INVX1 INVX1_687 ( .A(_5451_), .Y(_5626_) );
	AOI22X1 AOI22X1_844 ( .A(_5476_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_5626_), .Y(_5627_) );
	AOI22X1 AOI22X1_845 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_5550_), .C(_5429_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_5628_) );
	INVX1 INVX1_688 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_5629_) );
	INVX1 INVX1_689 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_5630_) );
	OAI22X1 OAI22X1_145 ( .A(_5629_), .B(_5438_), .C(_5436_), .D(_5630_), .Y(_5631_) );
	INVX1 INVX1_690 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_5632_) );
	NAND2X1 NAND2X1_1115 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_5539_), .Y(_5633_) );
	OAI21X1 OAI21X1_180 ( .A(_5632_), .B(_5444_), .C(_5633_), .Y(_5634_) );
	NOR2X1 NOR2X1_646 ( .A(_5631_), .B(_5634_), .Y(_5635_) );
	NAND3X1 NAND3X1_263 ( .A(_5627_), .B(_5628_), .C(_5635_), .Y(_5636_) );
	INVX1 INVX1_691 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_5637_) );
	NAND2X1 NAND2X1_1116 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_5423_), .Y(_5638_) );
	OAI21X1 OAI21X1_181 ( .A(_5637_), .B(_5453_), .C(_5638_), .Y(_5639_) );
	INVX1 INVX1_692 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_5640_) );
	INVX1 INVX1_693 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_5641_) );
	OAI22X1 OAI22X1_146 ( .A(_5640_), .B(_5459_), .C(_5457_), .D(_5641_), .Y(_5642_) );
	NOR2X1 NOR2X1_647 ( .A(_5642_), .B(_5639_), .Y(_5643_) );
	AOI22X1 AOI22X1_846 ( .A(_5543_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_5516_), .Y(_5644_) );
	AND2X2 AND2X2_117 ( .A(_5390_), .B(_5405_), .Y(_5645_) );
	AOI22X1 AOI22X1_847 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_5515_), .C(_5645_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_5646_) );
	NAND3X1 NAND3X1_264 ( .A(_5644_), .B(_5646_), .C(_5643_), .Y(_5647_) );
	NOR3X1 NOR3X1_470 ( .A(_5647_), .B(_5625_), .C(_5636_), .Y(_5648_) );
	INVX1 INVX1_694 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_5649_) );
	NAND2X1 NAND2X1_1117 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_5478_), .Y(_5650_) );
	OAI21X1 OAI21X1_182 ( .A(_5480_), .B(_5649_), .C(_5650_), .Y(_5651_) );
	AOI21X1 AOI21X1_128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_5527_), .C(_5651_), .Y(_5652_) );
	INVX1 INVX1_695 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_5653_) );
	INVX1 INVX1_696 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_5654_) );
	OAI22X1 OAI22X1_147 ( .A(_5654_), .B(_5486_), .C(_5487_), .D(_5653_), .Y(_5655_) );
	INVX1 INVX1_697 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_5656_) );
	NAND2X1 NAND2X1_1118 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_5496_), .Y(_5657_) );
	OAI21X1 OAI21X1_183 ( .A(_5397_), .B(_5656_), .C(_5657_), .Y(_5658_) );
	NOR2X1 NOR2X1_648 ( .A(_5658_), .B(_5655_), .Y(_5659_) );
	INVX1 INVX1_698 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_5660_) );
	INVX1 INVX1_699 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_5661_) );
	OAI22X1 OAI22X1_148 ( .A(_5492_), .B(_5661_), .C(_5498_), .D(_5660_), .Y(_5662_) );
	INVX1 INVX1_700 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_5663_) );
	NOR2X1 NOR2X1_649 ( .A(_5663_), .B(_5503_), .Y(_5664_) );
	INVX1 INVX1_701 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_5665_) );
	NOR2X1 NOR2X1_650 ( .A(_5665_), .B(_5504_), .Y(_5666_) );
	NOR3X1 NOR3X1_471 ( .A(_5664_), .B(_5662_), .C(_5666_), .Y(_5667_) );
	NAND3X1 NAND3X1_265 ( .A(_5659_), .B(_5652_), .C(_5667_), .Y(_5668_) );
	AOI22X1 AOI22X1_848 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_5508_), .C(_5509_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_5669_) );
	AOI22X1 AOI22X1_849 ( .A(_5511_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_5512_), .Y(_5670_) );
	NAND2X1 NAND2X1_1119 ( .A(_5669_), .B(_5670_), .Y(_5671_) );
	AOI22X1 AOI22X1_850 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_5519_), .C(_5518_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_5672_) );
	AOI22X1 AOI22X1_851 ( .A(_5462_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_5469_), .Y(_5673_) );
	NAND2X1 NAND2X1_1120 ( .A(_5672_), .B(_5673_), .Y(_5674_) );
	NOR2X1 NOR2X1_651 ( .A(_5671_), .B(_5674_), .Y(_5675_) );
	AOI22X1 AOI22X1_852 ( .A(_5523_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_5524_), .Y(_5676_) );
	AOI22X1 AOI22X1_853 ( .A(_5425_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_5526_), .Y(_5677_) );
	NAND2X1 NAND2X1_1121 ( .A(_5676_), .B(_5677_), .Y(_5678_) );
	AOI22X1 AOI22X1_854 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_5530_), .C(_5531_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_5679_) );
	AOI22X1 AOI22X1_855 ( .A(_5533_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_5534_), .Y(_5680_) );
	NAND2X1 NAND2X1_1122 ( .A(_5680_), .B(_5679_), .Y(_5681_) );
	NOR2X1 NOR2X1_652 ( .A(_5678_), .B(_5681_), .Y(_5682_) );
	NAND2X1 NAND2X1_1123 ( .A(_5682_), .B(_5675_), .Y(_5683_) );
	AOI22X1 AOI22X1_856 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_5540_), .C(_5441_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_5684_) );
	AOI22X1 AOI22X1_857 ( .A(_5464_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_5542_), .Y(_5685_) );
	NAND2X1 NAND2X1_1124 ( .A(_5684_), .B(_5685_), .Y(_5686_) );
	AOI22X1 AOI22X1_858 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_5431_), .C(_5551_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_5687_) );
	NAND2X1 NAND2X1_1125 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_5546_), .Y(_5688_) );
	NAND2X1 NAND2X1_1126 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_5548_), .Y(_5689_) );
	NAND3X1 NAND3X1_266 ( .A(_5688_), .B(_5689_), .C(_5687_), .Y(_5690_) );
	NOR2X1 NOR2X1_653 ( .A(_5690_), .B(_5686_), .Y(_5691_) );
	AOI22X1 AOI22X1_859 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_5555_), .C(_5556_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_5692_) );
	NAND2X1 NAND2X1_1127 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_5558_), .Y(_5693_) );
	NAND2X1 NAND2X1_1128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_5560_), .Y(_5694_) );
	NAND3X1 NAND3X1_267 ( .A(_5693_), .B(_5694_), .C(_5692_), .Y(_5695_) );
	AOI22X1 AOI22X1_860 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_5564_), .C(_5563_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_5696_) );
	AOI22X1 AOI22X1_861 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_5567_), .C(_5566_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_5697_) );
	NAND2X1 NAND2X1_1129 ( .A(_5696_), .B(_5697_), .Y(_5698_) );
	NOR2X1 NOR2X1_654 ( .A(_5698_), .B(_5695_), .Y(_5699_) );
	NAND2X1 NAND2X1_1130 ( .A(_5691_), .B(_5699_), .Y(_5700_) );
	NOR3X1 NOR3X1_472 ( .A(_5683_), .B(_5668_), .C(_5700_), .Y(_5701_) );
	AOI21X1 AOI21X1_129 ( .A(wData[21]), .B(_5577_), .C(_5382_), .Y(_5702_) );
	AOI22X1 AOI22X1_862 ( .A(_5580_), .B(wData[17]), .C(wData[1]), .D(_5608_), .Y(_5703_) );
	AOI22X1 AOI22X1_863 ( .A(_5601_), .B(wData[45]), .C(wData[25]), .D(_5584_), .Y(_5704_) );
	NAND3X1 NAND3X1_268 ( .A(_5702_), .B(_5704_), .C(_5703_), .Y(_5705_) );
	NAND3X1 NAND3X1_269 ( .A(wData[49]), .B(_5578_), .C(_5612_), .Y(_5706_) );
	AOI22X1 AOI22X1_864 ( .A(wData[61]), .B(_5600_), .C(_5588_), .D(wData[5]), .Y(_5707_) );
	AND2X2 AND2X2_118 ( .A(_5707_), .B(_5706_), .Y(_5708_) );
	AOI22X1 AOI22X1_865 ( .A(_5597_), .B(wData[57]), .C(wData[41]), .D(_5604_), .Y(_5709_) );
	AOI22X1 AOI22X1_866 ( .A(wData[53]), .B(_5598_), .C(_5594_), .D(wData[33]), .Y(_5710_) );
	AND2X2 AND2X2_119 ( .A(_5710_), .B(_5709_), .Y(_5711_) );
	AOI22X1 AOI22X1_867 ( .A(_5614_), .B(wData[9]), .C(wData[13]), .D(_5615_), .Y(_5712_) );
	AOI22X1 AOI22X1_868 ( .A(_5590_), .B(wData[29]), .C(wData[37]), .D(_5606_), .Y(_5713_) );
	AND2X2 AND2X2_120 ( .A(_5712_), .B(_5713_), .Y(_5714_) );
	NAND3X1 NAND3X1_270 ( .A(_5708_), .B(_5714_), .C(_5711_), .Y(_5715_) );
	NOR2X1 NOR2X1_655 ( .A(_5705_), .B(_5715_), .Y(_5716_) );
	AOI21X1 AOI21X1_130 ( .A(_5648_), .B(_5701_), .C(_5716_), .Y(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_1_) );
	AOI21X1 AOI21X1_131 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_5621_), .C(_5383_), .Y(_5717_) );
	INVX1 INVX1_702 ( .A(_5480_), .Y(_5718_) );
	AOI22X1 AOI22X1_869 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_5391_), .C(_5718_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_5719_) );
	INVX1 INVX1_703 ( .A(_5492_), .Y(_5720_) );
	AOI22X1 AOI22X1_870 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_5527_), .C(_5720_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_5721_) );
	NAND3X1 NAND3X1_271 ( .A(_5721_), .B(_5717_), .C(_5719_), .Y(_5722_) );
	AOI22X1 AOI22X1_871 ( .A(_5476_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_5626_), .Y(_5723_) );
	AOI22X1 AOI22X1_872 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_5425_), .C(_5398_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_5724_) );
	INVX1 INVX1_704 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_5725_) );
	NAND2X1 NAND2X1_1131 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_5515_), .Y(_5726_) );
	OAI21X1 OAI21X1_184 ( .A(_5725_), .B(_5487_), .C(_5726_), .Y(_5727_) );
	INVX1 INVX1_705 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_5728_) );
	NAND2X1 NAND2X1_1132 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_5441_), .Y(_5729_) );
	OAI21X1 OAI21X1_185 ( .A(_5728_), .B(_5444_), .C(_5729_), .Y(_5730_) );
	NOR2X1 NOR2X1_656 ( .A(_5727_), .B(_5730_), .Y(_5731_) );
	NAND3X1 NAND3X1_272 ( .A(_5723_), .B(_5724_), .C(_5731_), .Y(_5732_) );
	INVX1 INVX1_706 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_5733_) );
	NAND2X1 NAND2X1_1133 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_5423_), .Y(_5734_) );
	OAI21X1 OAI21X1_186 ( .A(_5733_), .B(_5453_), .C(_5734_), .Y(_5735_) );
	INVX1 INVX1_707 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_5736_) );
	INVX1 INVX1_708 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_5737_) );
	OAI22X1 OAI22X1_149 ( .A(_5736_), .B(_5459_), .C(_5457_), .D(_5737_), .Y(_5738_) );
	NOR2X1 NOR2X1_657 ( .A(_5738_), .B(_5735_), .Y(_5739_) );
	AOI22X1 AOI22X1_873 ( .A(_5543_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_5516_), .Y(_5740_) );
	AND2X2 AND2X2_121 ( .A(_5415_), .B(_5437_), .Y(_5741_) );
	AOI22X1 AOI22X1_874 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_5741_), .C(_5645_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_5742_) );
	NAND3X1 NAND3X1_273 ( .A(_5740_), .B(_5742_), .C(_5739_), .Y(_5743_) );
	NOR3X1 NOR3X1_473 ( .A(_5743_), .B(_5722_), .C(_5732_), .Y(_5744_) );
	INVX1 INVX1_709 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_5745_) );
	NOR3X1 NOR3X1_474 ( .A(_5745_), .B(_5410_), .C(_5409_), .Y(_5746_) );
	AND2X2 AND2X2_122 ( .A(_5431_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_5747_) );
	AND2X2 AND2X2_123 ( .A(_5551_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_5748_) );
	NOR3X1 NOR3X1_475 ( .A(_5748_), .B(_5747_), .C(_5746_), .Y(_5749_) );
	INVX1 INVX1_710 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_5750_) );
	INVX1 INVX1_711 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_5751_) );
	OAI22X1 OAI22X1_150 ( .A(_5751_), .B(_5486_), .C(_5436_), .D(_5750_), .Y(_5752_) );
	INVX1 INVX1_712 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_5753_) );
	INVX1 INVX1_713 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_5754_) );
	NAND2X1 NAND2X1_1134 ( .A(_5427_), .B(_5428_), .Y(_5755_) );
	OAI22X1 OAI22X1_151 ( .A(_5755_), .B(_5754_), .C(_5753_), .D(_5406_), .Y(_5756_) );
	NOR2X1 NOR2X1_658 ( .A(_5752_), .B(_5756_), .Y(_5757_) );
	INVX1 INVX1_714 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_5758_) );
	NOR3X1 NOR3X1_476 ( .A(_5387_), .B(_5404_), .C(_5395_), .Y(_5759_) );
	NAND2X1 NAND2X1_1135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_5759_), .Y(_5760_) );
	OAI21X1 OAI21X1_187 ( .A(_5416_), .B(_5758_), .C(_5760_), .Y(_5761_) );
	INVX1 INVX1_715 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_5762_) );
	INVX1 INVX1_716 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_5763_) );
	OAI22X1 OAI22X1_152 ( .A(_5503_), .B(_5763_), .C(_5762_), .D(_5504_), .Y(_5764_) );
	NOR2X1 NOR2X1_659 ( .A(_5761_), .B(_5764_), .Y(_5765_) );
	NAND3X1 NAND3X1_274 ( .A(_5749_), .B(_5765_), .C(_5757_), .Y(_5766_) );
	AOI22X1 AOI22X1_875 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_5508_), .C(_5509_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_5767_) );
	AOI22X1 AOI22X1_876 ( .A(_5511_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_5512_), .Y(_5768_) );
	NAND2X1 NAND2X1_1136 ( .A(_5767_), .B(_5768_), .Y(_5769_) );
	AOI22X1 AOI22X1_877 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_5519_), .C(_5518_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_5770_) );
	AOI22X1 AOI22X1_878 ( .A(_5462_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_5469_), .Y(_5771_) );
	NAND2X1 NAND2X1_1137 ( .A(_5770_), .B(_5771_), .Y(_5772_) );
	NOR2X1 NOR2X1_660 ( .A(_5769_), .B(_5772_), .Y(_5773_) );
	AOI22X1 AOI22X1_879 ( .A(_5523_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_5524_), .Y(_5774_) );
	AOI22X1 AOI22X1_880 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_5550_), .C(_5526_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_5775_) );
	NAND2X1 NAND2X1_1138 ( .A(_5775_), .B(_5774_), .Y(_5776_) );
	AOI22X1 AOI22X1_881 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_5530_), .C(_5531_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_5777_) );
	AOI22X1 AOI22X1_882 ( .A(_5533_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_5534_), .Y(_5778_) );
	NAND2X1 NAND2X1_1139 ( .A(_5778_), .B(_5777_), .Y(_5779_) );
	NOR2X1 NOR2X1_661 ( .A(_5776_), .B(_5779_), .Y(_5780_) );
	NAND2X1 NAND2X1_1140 ( .A(_5780_), .B(_5773_), .Y(_5781_) );
	AOI22X1 AOI22X1_883 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_5540_), .C(_5539_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_5782_) );
	AOI22X1 AOI22X1_884 ( .A(_5464_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_5542_), .Y(_5783_) );
	NAND2X1 NAND2X1_1141 ( .A(_5782_), .B(_5783_), .Y(_5784_) );
	AOI22X1 AOI22X1_885 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_5548_), .C(_5546_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_5785_) );
	AOI22X1 AOI22X1_886 ( .A(_5478_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_5496_), .Y(_5786_) );
	NAND2X1 NAND2X1_1142 ( .A(_5786_), .B(_5785_), .Y(_5787_) );
	NOR2X1 NOR2X1_662 ( .A(_5787_), .B(_5784_), .Y(_5788_) );
	AOI22X1 AOI22X1_887 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_5555_), .C(_5556_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_5789_) );
	NAND2X1 NAND2X1_1143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_5558_), .Y(_5790_) );
	NAND2X1 NAND2X1_1144 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_5560_), .Y(_5791_) );
	NAND3X1 NAND3X1_275 ( .A(_5790_), .B(_5791_), .C(_5789_), .Y(_5792_) );
	AOI22X1 AOI22X1_888 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_5564_), .C(_5563_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_5793_) );
	AOI22X1 AOI22X1_889 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_5567_), .C(_5566_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_5794_) );
	NAND2X1 NAND2X1_1145 ( .A(_5793_), .B(_5794_), .Y(_5795_) );
	NOR2X1 NOR2X1_663 ( .A(_5795_), .B(_5792_), .Y(_5796_) );
	NAND2X1 NAND2X1_1146 ( .A(_5788_), .B(_5796_), .Y(_5797_) );
	NOR3X1 NOR3X1_477 ( .A(_5781_), .B(_5766_), .C(_5797_), .Y(_5798_) );
	AOI22X1 AOI22X1_890 ( .A(_5604_), .B(wData[42]), .C(wData[38]), .D(_5606_), .Y(_5799_) );
	AOI22X1 AOI22X1_891 ( .A(_5601_), .B(wData[46]), .C(_5608_), .D(wData[2]), .Y(_5800_) );
	NAND2X1 NAND2X1_1147 ( .A(_5799_), .B(_5800_), .Y(_5801_) );
	AOI21X1 AOI21X1_132 ( .A(wData[34]), .B(_5594_), .C(_5801_), .Y(_5802_) );
	INVX1 INVX1_717 ( .A(wData[50]), .Y(_5803_) );
	AOI22X1 AOI22X1_892 ( .A(_5614_), .B(wData[10]), .C(wData[14]), .D(_5615_), .Y(_5804_) );
	OAI21X1 OAI21X1_188 ( .A(_5803_), .B(_5613_), .C(_5804_), .Y(_5805_) );
	AOI22X1 AOI22X1_893 ( .A(_5577_), .B(wData[22]), .C(wData[18]), .D(_5580_), .Y(_5806_) );
	NAND2X1 NAND2X1_1148 ( .A(wData[26]), .B(_5584_), .Y(_5807_) );
	AOI22X1 AOI22X1_894 ( .A(_5590_), .B(wData[30]), .C(wData[6]), .D(_5588_), .Y(_5808_) );
	NAND3X1 NAND3X1_276 ( .A(_5807_), .B(_5808_), .C(_5806_), .Y(_5809_) );
	NOR2X1 NOR2X1_664 ( .A(_5805_), .B(_5809_), .Y(_5810_) );
	NAND2X1 NAND2X1_1149 ( .A(wData[58]), .B(_5597_), .Y(_5811_) );
	NAND2X1 NAND2X1_1150 ( .A(wData[54]), .B(_5598_), .Y(_5812_) );
	NAND2X1 NAND2X1_1151 ( .A(_5811_), .B(_5812_), .Y(_5813_) );
	AOI21X1 AOI21X1_133 ( .A(wData[62]), .B(_5600_), .C(_5813_), .Y(_5814_) );
	NAND3X1 NAND3X1_277 ( .A(_5802_), .B(_5814_), .C(_5810_), .Y(_5815_) );
	NOR2X1 NOR2X1_665 ( .A(_5382_), .B(_5815_), .Y(_5816_) );
	AOI21X1 AOI21X1_134 ( .A(_5744_), .B(_5798_), .C(_5816_), .Y(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_2_) );
	AOI21X1 AOI21X1_135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_5626_), .C(_5383_), .Y(_5817_) );
	AOI22X1 AOI22X1_895 ( .A(_5398_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_5718_), .Y(_5818_) );
	AOI22X1 AOI22X1_896 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_5720_), .C(_5476_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_5819_) );
	NAND3X1 NAND3X1_278 ( .A(_5819_), .B(_5817_), .C(_5818_), .Y(_5820_) );
	AOI22X1 AOI22X1_897 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_5425_), .C(_5423_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_5821_) );
	AOI22X1 AOI22X1_898 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_5496_), .C(_5621_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_5822_) );
	INVX1 INVX1_718 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_5823_) );
	INVX1 INVX1_719 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_5824_) );
	OAI22X1 OAI22X1_153 ( .A(_5823_), .B(_5438_), .C(_5487_), .D(_5824_), .Y(_5825_) );
	INVX1 INVX1_720 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_5826_) );
	NAND2X1 NAND2X1_1152 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_5539_), .Y(_5827_) );
	OAI21X1 OAI21X1_189 ( .A(_5826_), .B(_5444_), .C(_5827_), .Y(_5828_) );
	NOR2X1 NOR2X1_666 ( .A(_5825_), .B(_5828_), .Y(_5829_) );
	NAND3X1 NAND3X1_279 ( .A(_5821_), .B(_5822_), .C(_5829_), .Y(_5830_) );
	AND2X2 AND2X2_124 ( .A(_5452_), .B(_5386_), .Y(_5831_) );
	AOI22X1 AOI22X1_899 ( .A(_5391_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_5831_), .Y(_5832_) );
	AND2X2 AND2X2_125 ( .A(_5450_), .B(_5415_), .Y(_5833_) );
	AND2X2 AND2X2_126 ( .A(_5458_), .B(_5415_), .Y(_5834_) );
	AOI22X1 AOI22X1_900 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_5834_), .C(_5833_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_5835_) );
	NAND2X1 NAND2X1_1153 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_5543_), .Y(_5836_) );
	NAND2X1 NAND2X1_1154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_5516_), .Y(_5837_) );
	NAND2X1 NAND2X1_1155 ( .A(_5836_), .B(_5837_), .Y(_5838_) );
	INVX1 INVX1_721 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_5839_) );
	NAND2X1 NAND2X1_1156 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_5515_), .Y(_5840_) );
	OAI21X1 OAI21X1_190 ( .A(_5839_), .B(_5468_), .C(_5840_), .Y(_5841_) );
	NOR2X1 NOR2X1_667 ( .A(_5838_), .B(_5841_), .Y(_5842_) );
	NAND3X1 NAND3X1_280 ( .A(_5832_), .B(_5835_), .C(_5842_), .Y(_5843_) );
	NOR3X1 NOR3X1_478 ( .A(_5830_), .B(_5820_), .C(_5843_), .Y(_5844_) );
	INVX1 INVX1_722 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_5845_) );
	NAND2X1 NAND2X1_1157 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_5431_), .Y(_5846_) );
	OAI21X1 OAI21X1_191 ( .A(_5436_), .B(_5845_), .C(_5846_), .Y(_5847_) );
	AOI21X1 AOI21X1_136 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_5411_), .C(_5847_), .Y(_5848_) );
	INVX1 INVX1_723 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_5849_) );
	INVX1 INVX1_724 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_5850_) );
	OAI22X1 OAI22X1_154 ( .A(_5755_), .B(_5850_), .C(_5849_), .D(_5406_), .Y(_5851_) );
	INVX1 INVX1_725 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_5852_) );
	NAND2X1 NAND2X1_1158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_5551_), .Y(_5853_) );
	OAI21X1 OAI21X1_192 ( .A(_5416_), .B(_5852_), .C(_5853_), .Y(_5854_) );
	NOR2X1 NOR2X1_668 ( .A(_5854_), .B(_5851_), .Y(_5855_) );
	INVX1 INVX1_726 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_5856_) );
	INVX1 INVX1_727 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_5857_) );
	OAI22X1 OAI22X1_155 ( .A(_5503_), .B(_5857_), .C(_5856_), .D(_5504_), .Y(_5858_) );
	INVX1 INVX1_728 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_5859_) );
	NAND2X1 NAND2X1_1159 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_5550_), .Y(_5860_) );
	OAI21X1 OAI21X1_193 ( .A(_5859_), .B(_5486_), .C(_5860_), .Y(_5861_) );
	NOR2X1 NOR2X1_669 ( .A(_5861_), .B(_5858_), .Y(_5862_) );
	NAND3X1 NAND3X1_281 ( .A(_5848_), .B(_5862_), .C(_5855_), .Y(_5863_) );
	AOI22X1 AOI22X1_901 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_5508_), .C(_5509_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_5864_) );
	AOI22X1 AOI22X1_902 ( .A(_5511_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_5512_), .Y(_5865_) );
	NAND2X1 NAND2X1_1160 ( .A(_5864_), .B(_5865_), .Y(_5866_) );
	AOI22X1 AOI22X1_903 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_5519_), .C(_5518_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_5867_) );
	AOI22X1 AOI22X1_904 ( .A(_5462_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_5469_), .Y(_5868_) );
	NAND2X1 NAND2X1_1161 ( .A(_5867_), .B(_5868_), .Y(_5869_) );
	NOR2X1 NOR2X1_670 ( .A(_5866_), .B(_5869_), .Y(_5870_) );
	AOI22X1 AOI22X1_905 ( .A(_5523_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_5524_), .Y(_5871_) );
	AOI22X1 AOI22X1_906 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_5759_), .C(_5526_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_5872_) );
	NAND2X1 NAND2X1_1162 ( .A(_5872_), .B(_5871_), .Y(_5873_) );
	AOI22X1 AOI22X1_907 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_5530_), .C(_5531_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_5874_) );
	AOI22X1 AOI22X1_908 ( .A(_5533_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_5534_), .Y(_5875_) );
	NAND2X1 NAND2X1_1163 ( .A(_5875_), .B(_5874_), .Y(_5876_) );
	NOR2X1 NOR2X1_671 ( .A(_5873_), .B(_5876_), .Y(_5877_) );
	NAND2X1 NAND2X1_1164 ( .A(_5877_), .B(_5870_), .Y(_5878_) );
	AOI22X1 AOI22X1_909 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_5540_), .C(_5441_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_5879_) );
	AOI22X1 AOI22X1_910 ( .A(_5464_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_5542_), .Y(_5880_) );
	NAND2X1 NAND2X1_1165 ( .A(_5879_), .B(_5880_), .Y(_5881_) );
	AOI22X1 AOI22X1_911 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_5548_), .C(_5546_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_5882_) );
	AOI22X1 AOI22X1_912 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_5478_), .C(_5527_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_5883_) );
	NAND2X1 NAND2X1_1166 ( .A(_5883_), .B(_5882_), .Y(_5884_) );
	NOR2X1 NOR2X1_672 ( .A(_5884_), .B(_5881_), .Y(_5885_) );
	AOI22X1 AOI22X1_913 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_5555_), .C(_5556_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_5886_) );
	NAND2X1 NAND2X1_1167 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_5558_), .Y(_5887_) );
	NAND2X1 NAND2X1_1168 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_5560_), .Y(_5888_) );
	NAND3X1 NAND3X1_282 ( .A(_5887_), .B(_5888_), .C(_5886_), .Y(_5889_) );
	AOI22X1 AOI22X1_914 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_5564_), .C(_5563_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_5890_) );
	AOI22X1 AOI22X1_915 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_5567_), .C(_5566_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_5891_) );
	NAND2X1 NAND2X1_1169 ( .A(_5890_), .B(_5891_), .Y(_5892_) );
	NOR2X1 NOR2X1_673 ( .A(_5892_), .B(_5889_), .Y(_5893_) );
	NAND2X1 NAND2X1_1170 ( .A(_5885_), .B(_5893_), .Y(_5894_) );
	NOR3X1 NOR3X1_479 ( .A(_5878_), .B(_5863_), .C(_5894_), .Y(_5895_) );
	NAND2X1 NAND2X1_1171 ( .A(wData[59]), .B(_5597_), .Y(_5896_) );
	OAI21X1 OAI21X1_194 ( .A(_5381_), .B(wBusy_bF_buf1), .C(_5896_), .Y(_5897_) );
	NAND2X1 NAND2X1_1172 ( .A(wData[7]), .B(_5588_), .Y(_5898_) );
	NAND2X1 NAND2X1_1173 ( .A(wData[55]), .B(_5598_), .Y(_5899_) );
	AOI22X1 AOI22X1_916 ( .A(wData[63]), .B(_5600_), .C(_5590_), .D(wData[31]), .Y(_5900_) );
	NAND3X1 NAND3X1_283 ( .A(_5898_), .B(_5899_), .C(_5900_), .Y(_5901_) );
	OR2X2 OR2X2_64 ( .A(_5901_), .B(_5897_), .Y(_5902_) );
	INVX1 INVX1_729 ( .A(wData[51]), .Y(_5903_) );
	NAND2X1 NAND2X1_1174 ( .A(wData[47]), .B(_5601_), .Y(_5904_) );
	OAI21X1 OAI21X1_195 ( .A(_5903_), .B(_5613_), .C(_5904_), .Y(_5905_) );
	AOI21X1 AOI21X1_137 ( .A(wData[3]), .B(_5608_), .C(_5905_), .Y(_5906_) );
	AOI22X1 AOI22X1_917 ( .A(_5614_), .B(wData[11]), .C(wData[15]), .D(_5615_), .Y(_5907_) );
	AOI22X1 AOI22X1_918 ( .A(_5577_), .B(wData[23]), .C(wData[27]), .D(_5584_), .Y(_5908_) );
	AND2X2 AND2X2_127 ( .A(_5907_), .B(_5908_), .Y(_5909_) );
	NAND2X1 NAND2X1_1175 ( .A(wData[39]), .B(_5606_), .Y(_5910_) );
	NAND2X1 NAND2X1_1176 ( .A(wData[43]), .B(_5604_), .Y(_5911_) );
	NAND2X1 NAND2X1_1177 ( .A(_5910_), .B(_5911_), .Y(_5912_) );
	NAND2X1 NAND2X1_1178 ( .A(wData[19]), .B(_5580_), .Y(_5913_) );
	NAND2X1 NAND2X1_1179 ( .A(wData[35]), .B(_5594_), .Y(_5914_) );
	NAND2X1 NAND2X1_1180 ( .A(_5913_), .B(_5914_), .Y(_5915_) );
	NOR2X1 NOR2X1_674 ( .A(_5912_), .B(_5915_), .Y(_5916_) );
	NAND3X1 NAND3X1_284 ( .A(_5909_), .B(_5906_), .C(_5916_), .Y(_5917_) );
	NOR2X1 NOR2X1_675 ( .A(_5902_), .B(_5917_), .Y(_5918_) );
	AOI21X1 AOI21X1_138 ( .A(_5844_), .B(_5895_), .C(_5918_), .Y(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_3_) );
	INVX1 INVX1_730 ( .A(wSelec[121]), .Y(_5919_) );
	NOR2X1 NOR2X1_676 ( .A(wBusy_bF_buf0), .B(_5919_), .Y(_5920_) );
	INVX1 INVX1_731 ( .A(_5920_), .Y(_5921_) );
	INVX1 INVX1_732 ( .A(wSelec[131]), .Y(_5922_) );
	NAND2X1 NAND2X1_1181 ( .A(wSelec[130]), .B(_5922_), .Y(_5923_) );
	INVX2 INVX2_19 ( .A(_5923_), .Y(_5924_) );
	OR2X2 OR2X2_65 ( .A(wSelec[127]), .B(wSelec[126]), .Y(_5925_) );
	INVX1 INVX1_733 ( .A(wSelec[129]), .Y(_5926_) );
	NAND2X1 NAND2X1_1182 ( .A(wSelec[128]), .B(_5926_), .Y(_5927_) );
	NOR2X1 NOR2X1_677 ( .A(_5925_), .B(_5927_), .Y(_5928_) );
	AND2X2 AND2X2_128 ( .A(_5928_), .B(_5924_), .Y(_5929_) );
	AOI21X1 AOI21X1_139 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_5929_), .C(_5921_), .Y(_5930_) );
	INVX1 INVX1_734 ( .A(wSelec[127]), .Y(_5931_) );
	NAND2X1 NAND2X1_1183 ( .A(wSelec[126]), .B(_5931_), .Y(_5932_) );
	OR2X2 OR2X2_66 ( .A(wSelec[128]), .B(wSelec[129]), .Y(_5933_) );
	NOR2X1 NOR2X1_678 ( .A(_5933_), .B(_5932_), .Y(_5934_) );
	NAND2X1 NAND2X1_1184 ( .A(_5924_), .B(_5934_), .Y(_5935_) );
	INVX1 INVX1_735 ( .A(_5935_), .Y(_5936_) );
	INVX1 INVX1_736 ( .A(wSelec[126]), .Y(_5937_) );
	NAND2X1 NAND2X1_1185 ( .A(wSelec[127]), .B(_5937_), .Y(_5938_) );
	INVX1 INVX1_737 ( .A(wSelec[128]), .Y(_5939_) );
	NAND2X1 NAND2X1_1186 ( .A(wSelec[129]), .B(_5939_), .Y(_5940_) );
	NOR2X1 NOR2X1_679 ( .A(_5938_), .B(_5940_), .Y(_5941_) );
	NAND2X1 NAND2X1_1187 ( .A(wSelec[130]), .B(wSelec[131]), .Y(_5942_) );
	INVX1 INVX1_738 ( .A(_5942_), .Y(_5943_) );
	NAND2X1 NAND2X1_1188 ( .A(_5943_), .B(_5941_), .Y(_5944_) );
	INVX1 INVX1_739 ( .A(_5944_), .Y(_5945_) );
	AOI22X1 AOI22X1_919 ( .A(_5936_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_5945_), .Y(_5946_) );
	OR2X2 OR2X2_67 ( .A(_5932_), .B(_5933_), .Y(_5947_) );
	OR2X2 OR2X2_68 ( .A(wSelec[130]), .B(wSelec[131]), .Y(_5948_) );
	NOR2X1 NOR2X1_680 ( .A(_5948_), .B(_5947_), .Y(_5949_) );
	NOR2X1 NOR2X1_681 ( .A(_5927_), .B(_5932_), .Y(_5950_) );
	INVX1 INVX1_740 ( .A(wSelec[130]), .Y(_5951_) );
	NAND2X1 NAND2X1_1189 ( .A(wSelec[131]), .B(_5951_), .Y(_5952_) );
	INVX2 INVX2_20 ( .A(_5952_), .Y(_5953_) );
	NAND2X1 NAND2X1_1190 ( .A(_5953_), .B(_5950_), .Y(_5954_) );
	INVX1 INVX1_741 ( .A(_5954_), .Y(_5955_) );
	AOI22X1 AOI22X1_920 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_5949_), .C(_5955_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_5956_) );
	NAND3X1 NAND3X1_285 ( .A(_5930_), .B(_5956_), .C(_5946_), .Y(_5957_) );
	NOR2X1 NOR2X1_682 ( .A(wSelec[127]), .B(wSelec[126]), .Y(_5958_) );
	NOR2X1 NOR2X1_683 ( .A(wSelec[128]), .B(wSelec[129]), .Y(_5959_) );
	NAND2X1 NAND2X1_1191 ( .A(_5958_), .B(_5959_), .Y(_5960_) );
	NOR2X1 NOR2X1_684 ( .A(_5923_), .B(_5960_), .Y(_5961_) );
	NAND2X1 NAND2X1_1192 ( .A(wSelec[127]), .B(wSelec[126]), .Y(_5962_) );
	NOR3X1 NOR3X1_480 ( .A(_5933_), .B(_5962_), .C(_5923_), .Y(_5963_) );
	AOI22X1 AOI22X1_921 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_5963_), .C(_5961_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_5964_) );
	INVX1 INVX1_742 ( .A(_5948_), .Y(_5965_) );
	NOR2X1 NOR2X1_685 ( .A(_5933_), .B(_5938_), .Y(_5966_) );
	AND2X2 AND2X2_129 ( .A(_5966_), .B(_5965_), .Y(_5967_) );
	NAND2X1 NAND2X1_1193 ( .A(wSelec[128]), .B(wSelec[129]), .Y(_5968_) );
	NOR3X1 NOR3X1_481 ( .A(_5942_), .B(_5962_), .C(_5968_), .Y(_5969_) );
	AOI22X1 AOI22X1_922 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_5969_), .C(_5967_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_5970_) );
	INVX1 INVX1_743 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_5971_) );
	INVX1 INVX1_744 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_5972_) );
	NOR2X1 NOR2X1_686 ( .A(_5932_), .B(_5940_), .Y(_5973_) );
	NAND2X1 NAND2X1_1194 ( .A(_5943_), .B(_5973_), .Y(_5974_) );
	NOR2X1 NOR2X1_687 ( .A(_5962_), .B(_5968_), .Y(_5975_) );
	NAND2X1 NAND2X1_1195 ( .A(_5975_), .B(_5953_), .Y(_5976_) );
	OAI22X1 OAI22X1_156 ( .A(_5971_), .B(_5976_), .C(_5974_), .D(_5972_), .Y(_5977_) );
	INVX1 INVX1_745 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_5978_) );
	NOR3X1 NOR3X1_482 ( .A(_5923_), .B(_5938_), .C(_5940_), .Y(_5979_) );
	NAND2X1 NAND2X1_1196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_5979_), .Y(_5980_) );
	NOR2X1 NOR2X1_688 ( .A(_5962_), .B(_5927_), .Y(_5981_) );
	NAND2X1 NAND2X1_1197 ( .A(_5953_), .B(_5981_), .Y(_5982_) );
	OAI21X1 OAI21X1_196 ( .A(_5978_), .B(_5982_), .C(_5980_), .Y(_5983_) );
	NOR2X1 NOR2X1_689 ( .A(_5977_), .B(_5983_), .Y(_5984_) );
	NAND3X1 NAND3X1_286 ( .A(_5964_), .B(_5970_), .C(_5984_), .Y(_5985_) );
	INVX1 INVX1_746 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_5986_) );
	INVX1 INVX1_747 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_5987_) );
	NOR2X1 NOR2X1_690 ( .A(_5927_), .B(_5938_), .Y(_5988_) );
	NAND2X1 NAND2X1_1198 ( .A(_5924_), .B(_5988_), .Y(_5989_) );
	NOR2X1 NOR2X1_691 ( .A(_5925_), .B(_5940_), .Y(_5990_) );
	NAND2X1 NAND2X1_1199 ( .A(_5924_), .B(_5990_), .Y(_5991_) );
	OAI22X1 OAI22X1_157 ( .A(_5991_), .B(_5986_), .C(_5987_), .D(_5989_), .Y(_5992_) );
	INVX1 INVX1_748 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_5993_) );
	INVX1 INVX1_749 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_5994_) );
	NAND2X1 NAND2X1_1200 ( .A(_5953_), .B(_5988_), .Y(_5995_) );
	NOR2X1 NOR2X1_692 ( .A(_5962_), .B(_5933_), .Y(_5996_) );
	NAND2X1 NAND2X1_1201 ( .A(_5953_), .B(_5996_), .Y(_5997_) );
	OAI22X1 OAI22X1_158 ( .A(_5993_), .B(_5997_), .C(_5995_), .D(_5994_), .Y(_5998_) );
	NOR2X1 NOR2X1_693 ( .A(_5998_), .B(_5992_), .Y(_5999_) );
	NOR3X1 NOR3X1_483 ( .A(_5932_), .B(_5968_), .C(_5952_), .Y(_6000_) );
	NAND2X1 NAND2X1_1202 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_6000_), .Y(_6001_) );
	NOR3X1 NOR3X1_484 ( .A(_5940_), .B(_5962_), .C(_5952_), .Y(_6002_) );
	NAND2X1 NAND2X1_1203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_6002_), .Y(_6003_) );
	NAND2X1 NAND2X1_1204 ( .A(_6001_), .B(_6003_), .Y(_6004_) );
	INVX1 INVX1_750 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_6005_) );
	NAND2X1 NAND2X1_1205 ( .A(_5943_), .B(_5928_), .Y(_6006_) );
	NOR3X1 NOR3X1_485 ( .A(_5938_), .B(_5940_), .C(_5952_), .Y(_6007_) );
	NAND2X1 NAND2X1_1206 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_6007_), .Y(_6008_) );
	OAI21X1 OAI21X1_197 ( .A(_6005_), .B(_6006_), .C(_6008_), .Y(_6009_) );
	NOR2X1 NOR2X1_694 ( .A(_6004_), .B(_6009_), .Y(_6010_) );
	NAND2X1 NAND2X1_1207 ( .A(_5999_), .B(_6010_), .Y(_6011_) );
	NOR3X1 NOR3X1_486 ( .A(_5957_), .B(_6011_), .C(_5985_), .Y(_6012_) );
	NAND2X1 NAND2X1_1208 ( .A(_5924_), .B(_5981_), .Y(_6013_) );
	INVX1 INVX1_751 ( .A(_6013_), .Y(_6014_) );
	INVX1 INVX1_752 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_6015_) );
	NOR3X1 NOR3X1_487 ( .A(_5925_), .B(_5948_), .C(_5927_), .Y(_6016_) );
	NAND2X1 NAND2X1_1209 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_6016_), .Y(_6017_) );
	NAND2X1 NAND2X1_1210 ( .A(_5965_), .B(_5988_), .Y(_6018_) );
	OAI21X1 OAI21X1_198 ( .A(_6018_), .B(_6015_), .C(_6017_), .Y(_6019_) );
	AOI21X1 AOI21X1_140 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_6014_), .C(_6019_), .Y(_6020_) );
	INVX1 INVX1_753 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_6021_) );
	INVX1 INVX1_754 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_6022_) );
	NOR2X1 NOR2X1_695 ( .A(_5968_), .B(_5925_), .Y(_6023_) );
	NAND2X1 NAND2X1_1211 ( .A(_5924_), .B(_6023_), .Y(_6024_) );
	NAND2X1 NAND2X1_1212 ( .A(_5965_), .B(_5950_), .Y(_6025_) );
	OAI22X1 OAI22X1_159 ( .A(_6022_), .B(_6024_), .C(_6025_), .D(_6021_), .Y(_6026_) );
	INVX1 INVX1_755 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_6027_) );
	INVX1 INVX1_756 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_6028_) );
	NAND2X1 NAND2X1_1213 ( .A(_5924_), .B(_5950_), .Y(_6029_) );
	NAND2X1 NAND2X1_1214 ( .A(_5965_), .B(_5996_), .Y(_6030_) );
	OAI22X1 OAI22X1_160 ( .A(_6027_), .B(_6030_), .C(_6029_), .D(_6028_), .Y(_6031_) );
	NOR2X1 NOR2X1_696 ( .A(_6026_), .B(_6031_), .Y(_6032_) );
	INVX1 INVX1_757 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_6033_) );
	NOR3X1 NOR3X1_488 ( .A(_5948_), .B(_5962_), .C(_5927_), .Y(_6034_) );
	NAND2X1 NAND2X1_1215 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_6034_), .Y(_6035_) );
	OR2X2 OR2X2_69 ( .A(_5960_), .B(_5942_), .Y(_6036_) );
	OAI21X1 OAI21X1_199 ( .A(_6033_), .B(_6036_), .C(_6035_), .Y(_6037_) );
	INVX1 INVX1_758 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_6038_) );
	INVX1 INVX1_759 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_6039_) );
	NOR2X1 NOR2X1_697 ( .A(_5968_), .B(_5938_), .Y(_6040_) );
	NAND2X1 NAND2X1_1216 ( .A(_5924_), .B(_6040_), .Y(_6041_) );
	NAND2X1 NAND2X1_1217 ( .A(_5943_), .B(_5934_), .Y(_6042_) );
	OAI22X1 OAI22X1_161 ( .A(_6041_), .B(_6039_), .C(_6038_), .D(_6042_), .Y(_6043_) );
	NOR2X1 NOR2X1_698 ( .A(_6037_), .B(_6043_), .Y(_6044_) );
	NAND3X1 NAND3X1_287 ( .A(_6020_), .B(_6044_), .C(_6032_), .Y(_6045_) );
	NOR3X1 NOR3X1_489 ( .A(_5925_), .B(_5933_), .C(_5948_), .Y(_6046_) );
	NOR3X1 NOR3X1_490 ( .A(_5942_), .B(_5968_), .C(_5932_), .Y(_6047_) );
	AOI22X1 AOI22X1_923 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_6046_), .C(_6047_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_6048_) );
	NOR3X1 NOR3X1_491 ( .A(_5942_), .B(_5968_), .C(_5938_), .Y(_6049_) );
	NOR3X1 NOR3X1_492 ( .A(_5942_), .B(_5962_), .C(_5940_), .Y(_6050_) );
	AOI22X1 AOI22X1_924 ( .A(_6049_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_6050_), .Y(_6051_) );
	NAND2X1 NAND2X1_1218 ( .A(_6048_), .B(_6051_), .Y(_6052_) );
	NOR3X1 NOR3X1_493 ( .A(_5940_), .B(_5925_), .C(_5952_), .Y(_6053_) );
	NOR3X1 NOR3X1_494 ( .A(_5932_), .B(_5940_), .C(_5952_), .Y(_6054_) );
	AOI22X1 AOI22X1_925 ( .A(_6053_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_6054_), .Y(_6055_) );
	NOR3X1 NOR3X1_495 ( .A(_5923_), .B(_5968_), .C(_5932_), .Y(_6056_) );
	NOR3X1 NOR3X1_496 ( .A(_5962_), .B(_5968_), .C(_5923_), .Y(_6057_) );
	AOI22X1 AOI22X1_926 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_6057_), .C(_6056_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_6058_) );
	NAND2X1 NAND2X1_1219 ( .A(_6058_), .B(_6055_), .Y(_6059_) );
	NOR2X1 NOR2X1_699 ( .A(_6052_), .B(_6059_), .Y(_6060_) );
	NOR3X1 NOR3X1_497 ( .A(_5948_), .B(_5968_), .C(_5932_), .Y(_6061_) );
	NOR3X1 NOR3X1_498 ( .A(_5948_), .B(_5968_), .C(_5938_), .Y(_6062_) );
	AOI22X1 AOI22X1_927 ( .A(_6061_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_6062_), .Y(_6063_) );
	NOR3X1 NOR3X1_499 ( .A(_5948_), .B(_5962_), .C(_5940_), .Y(_6064_) );
	NOR3X1 NOR3X1_500 ( .A(_5923_), .B(_5933_), .C(_5938_), .Y(_6065_) );
	AOI22X1 AOI22X1_928 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_6064_), .C(_6065_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_6066_) );
	NAND2X1 NAND2X1_1220 ( .A(_6063_), .B(_6066_), .Y(_6067_) );
	NOR3X1 NOR3X1_501 ( .A(_5962_), .B(_5968_), .C(_5948_), .Y(_6068_) );
	NOR3X1 NOR3X1_502 ( .A(_5938_), .B(_5933_), .C(_5952_), .Y(_6069_) );
	AOI22X1 AOI22X1_929 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_6068_), .C(_6069_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_6070_) );
	NOR3X1 NOR3X1_503 ( .A(_5925_), .B(_5933_), .C(_5952_), .Y(_6071_) );
	NOR3X1 NOR3X1_504 ( .A(_5925_), .B(_5968_), .C(_5952_), .Y(_6072_) );
	AOI22X1 AOI22X1_930 ( .A(_6071_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_6072_), .Y(_6073_) );
	NAND2X1 NAND2X1_1221 ( .A(_6073_), .B(_6070_), .Y(_6074_) );
	NOR2X1 NOR2X1_700 ( .A(_6067_), .B(_6074_), .Y(_6075_) );
	NAND2X1 NAND2X1_1222 ( .A(_6075_), .B(_6060_), .Y(_6076_) );
	NOR3X1 NOR3X1_505 ( .A(_5923_), .B(_5962_), .C(_5940_), .Y(_6077_) );
	NOR3X1 NOR3X1_506 ( .A(_5933_), .B(_5942_), .C(_5938_), .Y(_6078_) );
	AOI22X1 AOI22X1_931 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_6078_), .C(_6077_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_6079_) );
	NOR3X1 NOR3X1_507 ( .A(_5927_), .B(_5925_), .C(_5952_), .Y(_6080_) );
	NOR3X1 NOR3X1_508 ( .A(_5938_), .B(_5968_), .C(_5952_), .Y(_6081_) );
	AOI22X1 AOI22X1_932 ( .A(_6080_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_6081_), .Y(_6082_) );
	NAND2X1 NAND2X1_1223 ( .A(_6079_), .B(_6082_), .Y(_6083_) );
	NOR3X1 NOR3X1_509 ( .A(_5923_), .B(_5932_), .C(_5940_), .Y(_6084_) );
	NAND2X1 NAND2X1_1224 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_6084_), .Y(_6085_) );
	NOR3X1 NOR3X1_510 ( .A(_5942_), .B(_5962_), .C(_5927_), .Y(_6086_) );
	NAND2X1 NAND2X1_1225 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_6086_), .Y(_6087_) );
	NOR3X1 NOR3X1_511 ( .A(_5925_), .B(_5968_), .C(_5948_), .Y(_6088_) );
	NOR3X1 NOR3X1_512 ( .A(_5925_), .B(_5942_), .C(_5940_), .Y(_6089_) );
	AOI22X1 AOI22X1_933 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_6088_), .C(_6089_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_6090_) );
	NAND3X1 NAND3X1_288 ( .A(_6085_), .B(_6087_), .C(_6090_), .Y(_6091_) );
	NOR2X1 NOR2X1_701 ( .A(_6091_), .B(_6083_), .Y(_6092_) );
	NOR3X1 NOR3X1_513 ( .A(_5925_), .B(_5948_), .C(_5940_), .Y(_6093_) );
	NOR3X1 NOR3X1_514 ( .A(_5927_), .B(_5942_), .C(_5932_), .Y(_6094_) );
	AOI22X1 AOI22X1_934 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_6093_), .C(_6094_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_6095_) );
	NOR3X1 NOR3X1_515 ( .A(_5927_), .B(_5942_), .C(_5938_), .Y(_6096_) );
	NAND2X1 NAND2X1_1226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_6096_), .Y(_6097_) );
	NOR3X1 NOR3X1_516 ( .A(_5932_), .B(_5933_), .C(_5952_), .Y(_6098_) );
	NAND2X1 NAND2X1_1227 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_6098_), .Y(_6099_) );
	NAND3X1 NAND3X1_289 ( .A(_6097_), .B(_6099_), .C(_6095_), .Y(_6100_) );
	NOR3X1 NOR3X1_517 ( .A(_5932_), .B(_5948_), .C(_5940_), .Y(_6101_) );
	NOR3X1 NOR3X1_518 ( .A(_5942_), .B(_5968_), .C(_5925_), .Y(_6102_) );
	AOI22X1 AOI22X1_935 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_6102_), .C(_6101_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_6103_) );
	NOR3X1 NOR3X1_519 ( .A(_5938_), .B(_5948_), .C(_5940_), .Y(_6104_) );
	NOR3X1 NOR3X1_520 ( .A(_5942_), .B(_5962_), .C(_5933_), .Y(_6105_) );
	AOI22X1 AOI22X1_936 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_6105_), .C(_6104_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_6106_) );
	NAND2X1 NAND2X1_1228 ( .A(_6103_), .B(_6106_), .Y(_6107_) );
	NOR2X1 NOR2X1_702 ( .A(_6107_), .B(_6100_), .Y(_6108_) );
	NAND2X1 NAND2X1_1229 ( .A(_6092_), .B(_6108_), .Y(_6109_) );
	NOR3X1 NOR3X1_521 ( .A(_6076_), .B(_6045_), .C(_6109_), .Y(_6110_) );
	INVX1 INVX1_760 ( .A(wSelec[123]), .Y(_6111_) );
	NAND2X1 NAND2X1_1230 ( .A(wSelec[122]), .B(_6111_), .Y(_6112_) );
	INVX1 INVX1_761 ( .A(wSelec[125]), .Y(_6113_) );
	NAND2X1 NAND2X1_1231 ( .A(wSelec[124]), .B(_6113_), .Y(_6114_) );
	NOR2X1 NOR2X1_703 ( .A(_6112_), .B(_6114_), .Y(_6115_) );
	NOR2X1 NOR2X1_704 ( .A(wSelec[123]), .B(wSelec[122]), .Y(_6116_) );
	INVX1 INVX1_762 ( .A(_6116_), .Y(_6117_) );
	NOR2X1 NOR2X1_705 ( .A(_6114_), .B(_6117_), .Y(_6118_) );
	AOI22X1 AOI22X1_937 ( .A(wData[20]), .B(_6115_), .C(_6118_), .D(wData[16]), .Y(_6119_) );
	INVX1 INVX1_763 ( .A(wSelec[122]), .Y(_6120_) );
	NAND2X1 NAND2X1_1232 ( .A(wSelec[123]), .B(_6120_), .Y(_6121_) );
	NOR2X1 NOR2X1_706 ( .A(_6121_), .B(_6114_), .Y(_6122_) );
	NAND2X1 NAND2X1_1233 ( .A(wData[24]), .B(_6122_), .Y(_6123_) );
	INVX1 INVX1_764 ( .A(wSelec[124]), .Y(_6124_) );
	NAND2X1 NAND2X1_1234 ( .A(_6124_), .B(_6113_), .Y(_6125_) );
	NOR2X1 NOR2X1_707 ( .A(_6112_), .B(_6125_), .Y(_6126_) );
	NAND2X1 NAND2X1_1235 ( .A(wSelec[123]), .B(wSelec[122]), .Y(_6127_) );
	NOR2X1 NOR2X1_708 ( .A(_6127_), .B(_6114_), .Y(_6128_) );
	AOI22X1 AOI22X1_938 ( .A(_6128_), .B(wData[28]), .C(wData[4]), .D(_6126_), .Y(_6129_) );
	NAND3X1 NAND3X1_290 ( .A(_6123_), .B(_6129_), .C(_6119_), .Y(_6130_) );
	NAND2X1 NAND2X1_1236 ( .A(wSelec[125]), .B(_6124_), .Y(_6131_) );
	NOR2X1 NOR2X1_709 ( .A(_6131_), .B(_6117_), .Y(_6132_) );
	NAND2X1 NAND2X1_1237 ( .A(wData[32]), .B(_6132_), .Y(_6133_) );
	NAND2X1 NAND2X1_1238 ( .A(wSelec[124]), .B(wSelec[125]), .Y(_6134_) );
	NOR2X1 NOR2X1_710 ( .A(_6134_), .B(_6121_), .Y(_6135_) );
	NOR2X1 NOR2X1_711 ( .A(_6134_), .B(_6112_), .Y(_6136_) );
	AOI22X1 AOI22X1_939 ( .A(_6135_), .B(wData[56]), .C(wData[52]), .D(_6136_), .Y(_6137_) );
	NOR2X1 NOR2X1_712 ( .A(_6127_), .B(_6134_), .Y(_6138_) );
	NOR2X1 NOR2X1_713 ( .A(_6127_), .B(_6131_), .Y(_6139_) );
	AOI22X1 AOI22X1_940 ( .A(wData[60]), .B(_6138_), .C(_6139_), .D(wData[44]), .Y(_6140_) );
	NAND3X1 NAND3X1_291 ( .A(_6133_), .B(_6140_), .C(_6137_), .Y(_6141_) );
	NOR2X1 NOR2X1_714 ( .A(_6121_), .B(_6131_), .Y(_6142_) );
	NAND2X1 NAND2X1_1239 ( .A(wData[40]), .B(_6142_), .Y(_6143_) );
	NOR2X1 NOR2X1_715 ( .A(_6131_), .B(_6112_), .Y(_6144_) );
	NAND2X1 NAND2X1_1240 ( .A(wData[36]), .B(_6144_), .Y(_6145_) );
	NOR2X1 NOR2X1_716 ( .A(_6125_), .B(_6117_), .Y(_6146_) );
	NAND2X1 NAND2X1_1241 ( .A(wData[0]), .B(_6146_), .Y(_6147_) );
	NAND3X1 NAND3X1_292 ( .A(_6143_), .B(_6145_), .C(_6147_), .Y(_6148_) );
	INVX1 INVX1_765 ( .A(wData[48]), .Y(_6149_) );
	NOR2X1 NOR2X1_717 ( .A(_6124_), .B(_6113_), .Y(_6150_) );
	NAND2X1 NAND2X1_1242 ( .A(_6116_), .B(_6150_), .Y(_6151_) );
	NOR2X1 NOR2X1_718 ( .A(_6121_), .B(_6125_), .Y(_6152_) );
	NOR2X1 NOR2X1_719 ( .A(_6127_), .B(_6125_), .Y(_6153_) );
	AOI22X1 AOI22X1_941 ( .A(_6152_), .B(wData[8]), .C(wData[12]), .D(_6153_), .Y(_6154_) );
	OAI21X1 OAI21X1_200 ( .A(_6149_), .B(_6151_), .C(_6154_), .Y(_6155_) );
	OR2X2 OR2X2_70 ( .A(_6155_), .B(_6148_), .Y(_6156_) );
	NOR3X1 NOR3X1_522 ( .A(_6130_), .B(_6141_), .C(_6156_), .Y(_6157_) );
	AND2X2 AND2X2_130 ( .A(_6157_), .B(_5921_), .Y(_6158_) );
	AOI21X1 AOI21X1_141 ( .A(_6012_), .B(_6110_), .C(_6158_), .Y(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_0_) );
	INVX1 INVX1_766 ( .A(_6029_), .Y(_6159_) );
	AOI21X1 AOI21X1_142 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_6159_), .C(_5921_), .Y(_6160_) );
	AOI22X1 AOI22X1_942 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_5929_), .C(_5945_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_6161_) );
	AOI22X1 AOI22X1_943 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_5949_), .C(_5955_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_6162_) );
	NAND3X1 NAND3X1_293 ( .A(_6160_), .B(_6161_), .C(_6162_), .Y(_6163_) );
	INVX1 INVX1_767 ( .A(_5989_), .Y(_6164_) );
	AOI22X1 AOI22X1_944 ( .A(_6014_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_6164_), .Y(_6165_) );
	AOI22X1 AOI22X1_945 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_6088_), .C(_5967_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_6166_) );
	INVX1 INVX1_768 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_6167_) );
	INVX1 INVX1_769 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_6168_) );
	OAI22X1 OAI22X1_162 ( .A(_6167_), .B(_5976_), .C(_5974_), .D(_6168_), .Y(_6169_) );
	INVX1 INVX1_770 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_6170_) );
	NAND2X1 NAND2X1_1243 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_6077_), .Y(_6171_) );
	OAI21X1 OAI21X1_201 ( .A(_6170_), .B(_5982_), .C(_6171_), .Y(_6172_) );
	NOR2X1 NOR2X1_720 ( .A(_6169_), .B(_6172_), .Y(_6173_) );
	NAND3X1 NAND3X1_294 ( .A(_6165_), .B(_6166_), .C(_6173_), .Y(_6174_) );
	INVX1 INVX1_771 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_6175_) );
	NAND2X1 NAND2X1_1244 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_5961_), .Y(_6176_) );
	OAI21X1 OAI21X1_202 ( .A(_6175_), .B(_5991_), .C(_6176_), .Y(_6177_) );
	INVX1 INVX1_772 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_6178_) );
	INVX1 INVX1_773 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_6179_) );
	OAI22X1 OAI22X1_163 ( .A(_6178_), .B(_5997_), .C(_5995_), .D(_6179_), .Y(_6180_) );
	NOR2X1 NOR2X1_721 ( .A(_6180_), .B(_6177_), .Y(_6181_) );
	AOI22X1 AOI22X1_946 ( .A(_6081_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_6054_), .Y(_6182_) );
	AND2X2 AND2X2_131 ( .A(_5928_), .B(_5943_), .Y(_6183_) );
	AOI22X1 AOI22X1_947 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_6053_), .C(_6183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_6184_) );
	NAND3X1 NAND3X1_295 ( .A(_6182_), .B(_6184_), .C(_6181_), .Y(_6185_) );
	NOR3X1 NOR3X1_523 ( .A(_6185_), .B(_6163_), .C(_6174_), .Y(_6186_) );
	INVX1 INVX1_774 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_6187_) );
	NAND2X1 NAND2X1_1245 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_6016_), .Y(_6188_) );
	OAI21X1 OAI21X1_203 ( .A(_6018_), .B(_6187_), .C(_6188_), .Y(_6189_) );
	AOI21X1 AOI21X1_143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_6065_), .C(_6189_), .Y(_6190_) );
	INVX1 INVX1_775 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_6191_) );
	INVX1 INVX1_776 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_6192_) );
	OAI22X1 OAI22X1_164 ( .A(_6192_), .B(_6024_), .C(_6025_), .D(_6191_), .Y(_6193_) );
	INVX1 INVX1_777 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_6194_) );
	NAND2X1 NAND2X1_1246 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_6034_), .Y(_6195_) );
	OAI21X1 OAI21X1_204 ( .A(_5935_), .B(_6194_), .C(_6195_), .Y(_6196_) );
	NOR2X1 NOR2X1_722 ( .A(_6196_), .B(_6193_), .Y(_6197_) );
	INVX1 INVX1_778 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_6198_) );
	INVX1 INVX1_779 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_6199_) );
	OAI22X1 OAI22X1_165 ( .A(_6030_), .B(_6199_), .C(_6036_), .D(_6198_), .Y(_6200_) );
	INVX1 INVX1_780 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_6201_) );
	NOR2X1 NOR2X1_723 ( .A(_6201_), .B(_6041_), .Y(_6202_) );
	INVX1 INVX1_781 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_6203_) );
	NOR2X1 NOR2X1_724 ( .A(_6203_), .B(_6042_), .Y(_6204_) );
	NOR3X1 NOR3X1_524 ( .A(_6202_), .B(_6200_), .C(_6204_), .Y(_6205_) );
	NAND3X1 NAND3X1_296 ( .A(_6197_), .B(_6190_), .C(_6205_), .Y(_6206_) );
	AOI22X1 AOI22X1_948 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_6046_), .C(_6047_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_6207_) );
	AOI22X1 AOI22X1_949 ( .A(_6049_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_6050_), .Y(_6208_) );
	NAND2X1 NAND2X1_1247 ( .A(_6207_), .B(_6208_), .Y(_6209_) );
	AOI22X1 AOI22X1_950 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_6057_), .C(_6056_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_6210_) );
	AOI22X1 AOI22X1_951 ( .A(_6000_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_6007_), .Y(_6211_) );
	NAND2X1 NAND2X1_1248 ( .A(_6210_), .B(_6211_), .Y(_6212_) );
	NOR2X1 NOR2X1_725 ( .A(_6209_), .B(_6212_), .Y(_6213_) );
	AOI22X1 AOI22X1_952 ( .A(_6061_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_6062_), .Y(_6214_) );
	AOI22X1 AOI22X1_953 ( .A(_5963_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_6064_), .Y(_6215_) );
	NAND2X1 NAND2X1_1249 ( .A(_6214_), .B(_6215_), .Y(_6216_) );
	AOI22X1 AOI22X1_954 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_6068_), .C(_6069_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_6217_) );
	AOI22X1 AOI22X1_955 ( .A(_6071_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_6072_), .Y(_6218_) );
	NAND2X1 NAND2X1_1250 ( .A(_6218_), .B(_6217_), .Y(_6219_) );
	NOR2X1 NOR2X1_726 ( .A(_6216_), .B(_6219_), .Y(_6220_) );
	NAND2X1 NAND2X1_1251 ( .A(_6220_), .B(_6213_), .Y(_6221_) );
	AOI22X1 AOI22X1_956 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_6078_), .C(_5979_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_6222_) );
	AOI22X1 AOI22X1_957 ( .A(_6002_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_6080_), .Y(_6223_) );
	NAND2X1 NAND2X1_1252 ( .A(_6222_), .B(_6223_), .Y(_6224_) );
	AOI22X1 AOI22X1_958 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_5969_), .C(_6089_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_6225_) );
	NAND2X1 NAND2X1_1253 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_6084_), .Y(_6226_) );
	NAND2X1 NAND2X1_1254 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_6086_), .Y(_6227_) );
	NAND3X1 NAND3X1_297 ( .A(_6226_), .B(_6227_), .C(_6225_), .Y(_6228_) );
	NOR2X1 NOR2X1_727 ( .A(_6228_), .B(_6224_), .Y(_6229_) );
	AOI22X1 AOI22X1_959 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_6093_), .C(_6094_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_6230_) );
	NAND2X1 NAND2X1_1255 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_6096_), .Y(_6231_) );
	NAND2X1 NAND2X1_1256 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_6098_), .Y(_6232_) );
	NAND3X1 NAND3X1_298 ( .A(_6231_), .B(_6232_), .C(_6230_), .Y(_6233_) );
	AOI22X1 AOI22X1_960 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_6102_), .C(_6101_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_6234_) );
	AOI22X1 AOI22X1_961 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_6105_), .C(_6104_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_6235_) );
	NAND2X1 NAND2X1_1257 ( .A(_6234_), .B(_6235_), .Y(_6236_) );
	NOR2X1 NOR2X1_728 ( .A(_6236_), .B(_6233_), .Y(_6237_) );
	NAND2X1 NAND2X1_1258 ( .A(_6229_), .B(_6237_), .Y(_6238_) );
	NOR3X1 NOR3X1_525 ( .A(_6221_), .B(_6206_), .C(_6238_), .Y(_6239_) );
	AOI21X1 AOI21X1_144 ( .A(wData[21]), .B(_6115_), .C(_5920_), .Y(_6240_) );
	AOI22X1 AOI22X1_962 ( .A(_6118_), .B(wData[17]), .C(wData[1]), .D(_6146_), .Y(_6241_) );
	AOI22X1 AOI22X1_963 ( .A(_6139_), .B(wData[45]), .C(wData[25]), .D(_6122_), .Y(_6242_) );
	NAND3X1 NAND3X1_299 ( .A(_6240_), .B(_6242_), .C(_6241_), .Y(_6243_) );
	NAND3X1 NAND3X1_300 ( .A(wData[49]), .B(_6116_), .C(_6150_), .Y(_6244_) );
	AOI22X1 AOI22X1_964 ( .A(wData[61]), .B(_6138_), .C(_6126_), .D(wData[5]), .Y(_6245_) );
	AND2X2 AND2X2_132 ( .A(_6245_), .B(_6244_), .Y(_6246_) );
	AOI22X1 AOI22X1_965 ( .A(_6135_), .B(wData[57]), .C(wData[41]), .D(_6142_), .Y(_6247_) );
	AOI22X1 AOI22X1_966 ( .A(wData[53]), .B(_6136_), .C(_6132_), .D(wData[33]), .Y(_6248_) );
	AND2X2 AND2X2_133 ( .A(_6248_), .B(_6247_), .Y(_6249_) );
	AOI22X1 AOI22X1_967 ( .A(_6152_), .B(wData[9]), .C(wData[13]), .D(_6153_), .Y(_6250_) );
	AOI22X1 AOI22X1_968 ( .A(_6128_), .B(wData[29]), .C(wData[37]), .D(_6144_), .Y(_6251_) );
	AND2X2 AND2X2_134 ( .A(_6250_), .B(_6251_), .Y(_6252_) );
	NAND3X1 NAND3X1_301 ( .A(_6246_), .B(_6252_), .C(_6249_), .Y(_6253_) );
	NOR2X1 NOR2X1_729 ( .A(_6243_), .B(_6253_), .Y(_6254_) );
	AOI21X1 AOI21X1_145 ( .A(_6186_), .B(_6239_), .C(_6254_), .Y(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_1_) );
	AOI21X1 AOI21X1_146 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_6159_), .C(_5921_), .Y(_6255_) );
	INVX1 INVX1_782 ( .A(_6018_), .Y(_6256_) );
	AOI22X1 AOI22X1_969 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_5929_), .C(_6256_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_6257_) );
	INVX1 INVX1_783 ( .A(_6030_), .Y(_6258_) );
	AOI22X1 AOI22X1_970 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_6065_), .C(_6258_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_6259_) );
	NAND3X1 NAND3X1_302 ( .A(_6259_), .B(_6255_), .C(_6257_), .Y(_6260_) );
	AOI22X1 AOI22X1_971 ( .A(_6014_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_6164_), .Y(_6261_) );
	AOI22X1 AOI22X1_972 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_5963_), .C(_5936_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_6262_) );
	INVX1 INVX1_784 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_6263_) );
	NAND2X1 NAND2X1_1259 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_6053_), .Y(_6264_) );
	OAI21X1 OAI21X1_205 ( .A(_6263_), .B(_6025_), .C(_6264_), .Y(_6265_) );
	INVX1 INVX1_785 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_6266_) );
	NAND2X1 NAND2X1_1260 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_5979_), .Y(_6267_) );
	OAI21X1 OAI21X1_206 ( .A(_6266_), .B(_5982_), .C(_6267_), .Y(_6268_) );
	NOR2X1 NOR2X1_730 ( .A(_6265_), .B(_6268_), .Y(_6269_) );
	NAND3X1 NAND3X1_303 ( .A(_6261_), .B(_6262_), .C(_6269_), .Y(_6270_) );
	INVX1 INVX1_786 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_6271_) );
	NAND2X1 NAND2X1_1261 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_5961_), .Y(_6272_) );
	OAI21X1 OAI21X1_207 ( .A(_6271_), .B(_5991_), .C(_6272_), .Y(_6273_) );
	INVX1 INVX1_787 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_6274_) );
	INVX1 INVX1_788 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_6275_) );
	OAI22X1 OAI22X1_166 ( .A(_6274_), .B(_5997_), .C(_5995_), .D(_6275_), .Y(_6276_) );
	NOR2X1 NOR2X1_731 ( .A(_6276_), .B(_6273_), .Y(_6277_) );
	AOI22X1 AOI22X1_973 ( .A(_6081_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_6054_), .Y(_6278_) );
	AND2X2 AND2X2_135 ( .A(_5953_), .B(_5975_), .Y(_6279_) );
	AOI22X1 AOI22X1_974 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_6279_), .C(_6183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_6280_) );
	NAND3X1 NAND3X1_304 ( .A(_6278_), .B(_6280_), .C(_6277_), .Y(_6281_) );
	NOR3X1 NOR3X1_526 ( .A(_6281_), .B(_6260_), .C(_6270_), .Y(_6282_) );
	INVX1 INVX1_789 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_6283_) );
	NOR3X1 NOR3X1_527 ( .A(_6283_), .B(_5948_), .C(_5947_), .Y(_6284_) );
	AND2X2 AND2X2_136 ( .A(_5969_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_6285_) );
	AND2X2 AND2X2_137 ( .A(_6089_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_6286_) );
	NOR3X1 NOR3X1_528 ( .A(_6286_), .B(_6285_), .C(_6284_), .Y(_6287_) );
	INVX1 INVX1_790 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_6288_) );
	INVX1 INVX1_791 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_6289_) );
	OAI22X1 OAI22X1_167 ( .A(_6289_), .B(_6024_), .C(_5974_), .D(_6288_), .Y(_6290_) );
	INVX1 INVX1_792 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_6291_) );
	INVX1 INVX1_793 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_6292_) );
	NAND2X1 NAND2X1_1262 ( .A(_5965_), .B(_5966_), .Y(_6293_) );
	OAI22X1 OAI22X1_168 ( .A(_6293_), .B(_6292_), .C(_6291_), .D(_5944_), .Y(_6294_) );
	NOR2X1 NOR2X1_732 ( .A(_6290_), .B(_6294_), .Y(_6295_) );
	INVX1 INVX1_794 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_6296_) );
	NOR3X1 NOR3X1_529 ( .A(_5925_), .B(_5942_), .C(_5933_), .Y(_6297_) );
	NAND2X1 NAND2X1_1263 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_6297_), .Y(_6298_) );
	OAI21X1 OAI21X1_208 ( .A(_5954_), .B(_6296_), .C(_6298_), .Y(_6299_) );
	INVX1 INVX1_795 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_6300_) );
	INVX1 INVX1_796 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_6301_) );
	OAI22X1 OAI22X1_169 ( .A(_6041_), .B(_6301_), .C(_6300_), .D(_6042_), .Y(_6302_) );
	NOR2X1 NOR2X1_733 ( .A(_6299_), .B(_6302_), .Y(_6303_) );
	NAND3X1 NAND3X1_305 ( .A(_6287_), .B(_6303_), .C(_6295_), .Y(_6304_) );
	AOI22X1 AOI22X1_975 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_6046_), .C(_6047_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_6305_) );
	AOI22X1 AOI22X1_976 ( .A(_6049_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_6050_), .Y(_6306_) );
	NAND2X1 NAND2X1_1264 ( .A(_6305_), .B(_6306_), .Y(_6307_) );
	AOI22X1 AOI22X1_977 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_6057_), .C(_6056_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_6308_) );
	AOI22X1 AOI22X1_978 ( .A(_6000_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_6007_), .Y(_6309_) );
	NAND2X1 NAND2X1_1265 ( .A(_6308_), .B(_6309_), .Y(_6310_) );
	NOR2X1 NOR2X1_734 ( .A(_6307_), .B(_6310_), .Y(_6311_) );
	AOI22X1 AOI22X1_979 ( .A(_6061_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_6062_), .Y(_6312_) );
	AOI22X1 AOI22X1_980 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_6088_), .C(_6064_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_6313_) );
	NAND2X1 NAND2X1_1266 ( .A(_6313_), .B(_6312_), .Y(_6314_) );
	AOI22X1 AOI22X1_981 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_6068_), .C(_6069_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_6315_) );
	AOI22X1 AOI22X1_982 ( .A(_6071_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_6072_), .Y(_6316_) );
	NAND2X1 NAND2X1_1267 ( .A(_6316_), .B(_6315_), .Y(_6317_) );
	NOR2X1 NOR2X1_735 ( .A(_6314_), .B(_6317_), .Y(_6318_) );
	NAND2X1 NAND2X1_1268 ( .A(_6318_), .B(_6311_), .Y(_6319_) );
	AOI22X1 AOI22X1_983 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_6078_), .C(_6077_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_6320_) );
	AOI22X1 AOI22X1_984 ( .A(_6002_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_6080_), .Y(_6321_) );
	NAND2X1 NAND2X1_1269 ( .A(_6320_), .B(_6321_), .Y(_6322_) );
	AOI22X1 AOI22X1_985 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_6086_), .C(_6084_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_6323_) );
	AOI22X1 AOI22X1_986 ( .A(_6016_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_6034_), .Y(_6324_) );
	NAND2X1 NAND2X1_1270 ( .A(_6324_), .B(_6323_), .Y(_6325_) );
	NOR2X1 NOR2X1_736 ( .A(_6325_), .B(_6322_), .Y(_6326_) );
	AOI22X1 AOI22X1_987 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_6093_), .C(_6094_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_6327_) );
	NAND2X1 NAND2X1_1271 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_6096_), .Y(_6328_) );
	NAND2X1 NAND2X1_1272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_6098_), .Y(_6329_) );
	NAND3X1 NAND3X1_306 ( .A(_6328_), .B(_6329_), .C(_6327_), .Y(_6330_) );
	AOI22X1 AOI22X1_988 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_6102_), .C(_6101_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_6331_) );
	AOI22X1 AOI22X1_989 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_6105_), .C(_6104_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_6332_) );
	NAND2X1 NAND2X1_1273 ( .A(_6331_), .B(_6332_), .Y(_6333_) );
	NOR2X1 NOR2X1_737 ( .A(_6333_), .B(_6330_), .Y(_6334_) );
	NAND2X1 NAND2X1_1274 ( .A(_6326_), .B(_6334_), .Y(_6335_) );
	NOR3X1 NOR3X1_530 ( .A(_6319_), .B(_6304_), .C(_6335_), .Y(_6336_) );
	AOI22X1 AOI22X1_990 ( .A(_6142_), .B(wData[42]), .C(wData[38]), .D(_6144_), .Y(_6337_) );
	AOI22X1 AOI22X1_991 ( .A(_6139_), .B(wData[46]), .C(_6146_), .D(wData[2]), .Y(_6338_) );
	NAND2X1 NAND2X1_1275 ( .A(_6337_), .B(_6338_), .Y(_6339_) );
	AOI21X1 AOI21X1_147 ( .A(wData[34]), .B(_6132_), .C(_6339_), .Y(_6340_) );
	INVX1 INVX1_797 ( .A(wData[50]), .Y(_6341_) );
	AOI22X1 AOI22X1_992 ( .A(_6152_), .B(wData[10]), .C(wData[14]), .D(_6153_), .Y(_6342_) );
	OAI21X1 OAI21X1_209 ( .A(_6341_), .B(_6151_), .C(_6342_), .Y(_6343_) );
	AOI22X1 AOI22X1_993 ( .A(_6115_), .B(wData[22]), .C(wData[18]), .D(_6118_), .Y(_6344_) );
	NAND2X1 NAND2X1_1276 ( .A(wData[26]), .B(_6122_), .Y(_6345_) );
	AOI22X1 AOI22X1_994 ( .A(_6128_), .B(wData[30]), .C(wData[6]), .D(_6126_), .Y(_6346_) );
	NAND3X1 NAND3X1_307 ( .A(_6345_), .B(_6346_), .C(_6344_), .Y(_6347_) );
	NOR2X1 NOR2X1_738 ( .A(_6343_), .B(_6347_), .Y(_6348_) );
	NAND2X1 NAND2X1_1277 ( .A(wData[58]), .B(_6135_), .Y(_6349_) );
	NAND2X1 NAND2X1_1278 ( .A(wData[54]), .B(_6136_), .Y(_6350_) );
	NAND2X1 NAND2X1_1279 ( .A(_6349_), .B(_6350_), .Y(_6351_) );
	AOI21X1 AOI21X1_148 ( .A(wData[62]), .B(_6138_), .C(_6351_), .Y(_6352_) );
	NAND3X1 NAND3X1_308 ( .A(_6340_), .B(_6352_), .C(_6348_), .Y(_6353_) );
	NOR2X1 NOR2X1_739 ( .A(_5920_), .B(_6353_), .Y(_6354_) );
	AOI21X1 AOI21X1_149 ( .A(_6282_), .B(_6336_), .C(_6354_), .Y(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_2_) );
	AOI21X1 AOI21X1_150 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_6164_), .C(_5921_), .Y(_6355_) );
	AOI22X1 AOI22X1_995 ( .A(_5936_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_6256_), .Y(_6356_) );
	AOI22X1 AOI22X1_996 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_6258_), .C(_6014_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_6357_) );
	NAND3X1 NAND3X1_309 ( .A(_6357_), .B(_6355_), .C(_6356_), .Y(_6358_) );
	AOI22X1 AOI22X1_997 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_5963_), .C(_5961_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_6359_) );
	AOI22X1 AOI22X1_998 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_6034_), .C(_6159_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_6360_) );
	INVX1 INVX1_798 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_6361_) );
	INVX1 INVX1_799 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_6362_) );
	OAI22X1 OAI22X1_170 ( .A(_6361_), .B(_5976_), .C(_6025_), .D(_6362_), .Y(_6363_) );
	INVX1 INVX1_800 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_6364_) );
	NAND2X1 NAND2X1_1280 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_6077_), .Y(_6365_) );
	OAI21X1 OAI21X1_210 ( .A(_6364_), .B(_5982_), .C(_6365_), .Y(_6366_) );
	NOR2X1 NOR2X1_740 ( .A(_6363_), .B(_6366_), .Y(_6367_) );
	NAND3X1 NAND3X1_310 ( .A(_6359_), .B(_6360_), .C(_6367_), .Y(_6368_) );
	AND2X2 AND2X2_138 ( .A(_5990_), .B(_5924_), .Y(_6369_) );
	AOI22X1 AOI22X1_999 ( .A(_5929_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_6369_), .Y(_6370_) );
	AND2X2 AND2X2_139 ( .A(_5988_), .B(_5953_), .Y(_6371_) );
	AND2X2 AND2X2_140 ( .A(_5996_), .B(_5953_), .Y(_6372_) );
	AOI22X1 AOI22X1_1000 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_6372_), .C(_6371_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_6373_) );
	NAND2X1 NAND2X1_1281 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_6081_), .Y(_6374_) );
	NAND2X1 NAND2X1_1282 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_6054_), .Y(_6375_) );
	NAND2X1 NAND2X1_1283 ( .A(_6374_), .B(_6375_), .Y(_6376_) );
	INVX1 INVX1_801 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_6377_) );
	NAND2X1 NAND2X1_1284 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_6053_), .Y(_6378_) );
	OAI21X1 OAI21X1_211 ( .A(_6377_), .B(_6006_), .C(_6378_), .Y(_6379_) );
	NOR2X1 NOR2X1_741 ( .A(_6376_), .B(_6379_), .Y(_6380_) );
	NAND3X1 NAND3X1_311 ( .A(_6370_), .B(_6373_), .C(_6380_), .Y(_6381_) );
	NOR3X1 NOR3X1_531 ( .A(_6368_), .B(_6358_), .C(_6381_), .Y(_6382_) );
	INVX1 INVX1_802 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_6383_) );
	NAND2X1 NAND2X1_1285 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_5969_), .Y(_6384_) );
	OAI21X1 OAI21X1_212 ( .A(_5974_), .B(_6383_), .C(_6384_), .Y(_6385_) );
	AOI21X1 AOI21X1_151 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_5949_), .C(_6385_), .Y(_6386_) );
	INVX1 INVX1_803 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_6387_) );
	INVX1 INVX1_804 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_6388_) );
	OAI22X1 OAI22X1_171 ( .A(_6293_), .B(_6388_), .C(_6387_), .D(_5944_), .Y(_6389_) );
	INVX1 INVX1_805 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_6390_) );
	NAND2X1 NAND2X1_1286 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_6089_), .Y(_6391_) );
	OAI21X1 OAI21X1_213 ( .A(_5954_), .B(_6390_), .C(_6391_), .Y(_6392_) );
	NOR2X1 NOR2X1_742 ( .A(_6392_), .B(_6389_), .Y(_6393_) );
	INVX1 INVX1_806 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_6394_) );
	INVX1 INVX1_807 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_6395_) );
	OAI22X1 OAI22X1_172 ( .A(_6041_), .B(_6395_), .C(_6394_), .D(_6042_), .Y(_6396_) );
	INVX1 INVX1_808 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_6397_) );
	NAND2X1 NAND2X1_1287 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_6088_), .Y(_6398_) );
	OAI21X1 OAI21X1_214 ( .A(_6397_), .B(_6024_), .C(_6398_), .Y(_6399_) );
	NOR2X1 NOR2X1_743 ( .A(_6399_), .B(_6396_), .Y(_6400_) );
	NAND3X1 NAND3X1_312 ( .A(_6386_), .B(_6400_), .C(_6393_), .Y(_6401_) );
	AOI22X1 AOI22X1_1001 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_6046_), .C(_6047_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_6402_) );
	AOI22X1 AOI22X1_1002 ( .A(_6049_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_6050_), .Y(_6403_) );
	NAND2X1 NAND2X1_1288 ( .A(_6402_), .B(_6403_), .Y(_6404_) );
	AOI22X1 AOI22X1_1003 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_6057_), .C(_6056_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_6405_) );
	AOI22X1 AOI22X1_1004 ( .A(_6000_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_6007_), .Y(_6406_) );
	NAND2X1 NAND2X1_1289 ( .A(_6405_), .B(_6406_), .Y(_6407_) );
	NOR2X1 NOR2X1_744 ( .A(_6404_), .B(_6407_), .Y(_6408_) );
	AOI22X1 AOI22X1_1005 ( .A(_6061_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_6062_), .Y(_6409_) );
	AOI22X1 AOI22X1_1006 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_6297_), .C(_6064_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_6410_) );
	NAND2X1 NAND2X1_1290 ( .A(_6410_), .B(_6409_), .Y(_6411_) );
	AOI22X1 AOI22X1_1007 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_6068_), .C(_6069_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_6412_) );
	AOI22X1 AOI22X1_1008 ( .A(_6071_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_6072_), .Y(_6413_) );
	NAND2X1 NAND2X1_1291 ( .A(_6413_), .B(_6412_), .Y(_6414_) );
	NOR2X1 NOR2X1_745 ( .A(_6411_), .B(_6414_), .Y(_6415_) );
	NAND2X1 NAND2X1_1292 ( .A(_6415_), .B(_6408_), .Y(_6416_) );
	AOI22X1 AOI22X1_1009 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_6078_), .C(_5979_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_6417_) );
	AOI22X1 AOI22X1_1010 ( .A(_6002_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_6080_), .Y(_6418_) );
	NAND2X1 NAND2X1_1293 ( .A(_6417_), .B(_6418_), .Y(_6419_) );
	AOI22X1 AOI22X1_1011 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_6086_), .C(_6084_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_6420_) );
	AOI22X1 AOI22X1_1012 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_6016_), .C(_6065_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_6421_) );
	NAND2X1 NAND2X1_1294 ( .A(_6421_), .B(_6420_), .Y(_6422_) );
	NOR2X1 NOR2X1_746 ( .A(_6422_), .B(_6419_), .Y(_6423_) );
	AOI22X1 AOI22X1_1013 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_6093_), .C(_6094_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_6424_) );
	NAND2X1 NAND2X1_1295 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_6096_), .Y(_6425_) );
	NAND2X1 NAND2X1_1296 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_6098_), .Y(_6426_) );
	NAND3X1 NAND3X1_313 ( .A(_6425_), .B(_6426_), .C(_6424_), .Y(_6427_) );
	AOI22X1 AOI22X1_1014 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_6102_), .C(_6101_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_6428_) );
	AOI22X1 AOI22X1_1015 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_6105_), .C(_6104_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_6429_) );
	NAND2X1 NAND2X1_1297 ( .A(_6428_), .B(_6429_), .Y(_6430_) );
	NOR2X1 NOR2X1_747 ( .A(_6430_), .B(_6427_), .Y(_6431_) );
	NAND2X1 NAND2X1_1298 ( .A(_6423_), .B(_6431_), .Y(_6432_) );
	NOR3X1 NOR3X1_532 ( .A(_6416_), .B(_6401_), .C(_6432_), .Y(_6433_) );
	NAND2X1 NAND2X1_1299 ( .A(wData[59]), .B(_6135_), .Y(_6434_) );
	OAI21X1 OAI21X1_215 ( .A(_5919_), .B(wBusy_bF_buf4), .C(_6434_), .Y(_6435_) );
	NAND2X1 NAND2X1_1300 ( .A(wData[7]), .B(_6126_), .Y(_6436_) );
	NAND2X1 NAND2X1_1301 ( .A(wData[55]), .B(_6136_), .Y(_6437_) );
	AOI22X1 AOI22X1_1016 ( .A(wData[63]), .B(_6138_), .C(_6128_), .D(wData[31]), .Y(_6438_) );
	NAND3X1 NAND3X1_314 ( .A(_6436_), .B(_6437_), .C(_6438_), .Y(_6439_) );
	OR2X2 OR2X2_71 ( .A(_6439_), .B(_6435_), .Y(_6440_) );
	INVX1 INVX1_809 ( .A(wData[51]), .Y(_6441_) );
	NAND2X1 NAND2X1_1302 ( .A(wData[47]), .B(_6139_), .Y(_6442_) );
	OAI21X1 OAI21X1_216 ( .A(_6441_), .B(_6151_), .C(_6442_), .Y(_6443_) );
	AOI21X1 AOI21X1_152 ( .A(wData[3]), .B(_6146_), .C(_6443_), .Y(_6444_) );
	AOI22X1 AOI22X1_1017 ( .A(_6152_), .B(wData[11]), .C(wData[15]), .D(_6153_), .Y(_6445_) );
	AOI22X1 AOI22X1_1018 ( .A(_6115_), .B(wData[23]), .C(wData[27]), .D(_6122_), .Y(_6446_) );
	AND2X2 AND2X2_141 ( .A(_6445_), .B(_6446_), .Y(_6447_) );
	NAND2X1 NAND2X1_1303 ( .A(wData[39]), .B(_6144_), .Y(_6448_) );
	NAND2X1 NAND2X1_1304 ( .A(wData[43]), .B(_6142_), .Y(_6449_) );
	NAND2X1 NAND2X1_1305 ( .A(_6448_), .B(_6449_), .Y(_6450_) );
	NAND2X1 NAND2X1_1306 ( .A(wData[19]), .B(_6118_), .Y(_6451_) );
	NAND2X1 NAND2X1_1307 ( .A(wData[35]), .B(_6132_), .Y(_6452_) );
	NAND2X1 NAND2X1_1308 ( .A(_6451_), .B(_6452_), .Y(_6453_) );
	NOR2X1 NOR2X1_748 ( .A(_6450_), .B(_6453_), .Y(_6454_) );
	NAND3X1 NAND3X1_315 ( .A(_6447_), .B(_6444_), .C(_6454_), .Y(_6455_) );
	NOR2X1 NOR2X1_749 ( .A(_6440_), .B(_6455_), .Y(_6456_) );
	AOI21X1 AOI21X1_153 ( .A(_6382_), .B(_6433_), .C(_6456_), .Y(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_3_) );
	INVX1 INVX1_810 ( .A(wSelec[132]), .Y(_6457_) );
	NOR2X1 NOR2X1_750 ( .A(wBusy_bF_buf3), .B(_6457_), .Y(_6458_) );
	INVX1 INVX1_811 ( .A(_6458_), .Y(_6459_) );
	INVX1 INVX1_812 ( .A(wSelec[142]), .Y(_6460_) );
	NAND2X1 NAND2X1_1309 ( .A(wSelec[141]), .B(_6460_), .Y(_6461_) );
	INVX2 INVX2_21 ( .A(_6461_), .Y(_6462_) );
	OR2X2 OR2X2_72 ( .A(wSelec[138]), .B(wSelec[137]), .Y(_6463_) );
	INVX1 INVX1_813 ( .A(wSelec[140]), .Y(_6464_) );
	NAND2X1 NAND2X1_1310 ( .A(wSelec[139]), .B(_6464_), .Y(_6465_) );
	NOR2X1 NOR2X1_751 ( .A(_6463_), .B(_6465_), .Y(_6466_) );
	AND2X2 AND2X2_142 ( .A(_6466_), .B(_6462_), .Y(_6467_) );
	AOI21X1 AOI21X1_154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_6467_), .C(_6459_), .Y(_6468_) );
	INVX1 INVX1_814 ( .A(wSelec[138]), .Y(_6469_) );
	NAND2X1 NAND2X1_1311 ( .A(wSelec[137]), .B(_6469_), .Y(_6470_) );
	OR2X2 OR2X2_73 ( .A(wSelec[139]), .B(wSelec[140]), .Y(_6471_) );
	NOR2X1 NOR2X1_752 ( .A(_6471_), .B(_6470_), .Y(_6472_) );
	NAND2X1 NAND2X1_1312 ( .A(_6462_), .B(_6472_), .Y(_6473_) );
	INVX1 INVX1_815 ( .A(_6473_), .Y(_6474_) );
	INVX1 INVX1_816 ( .A(wSelec[137]), .Y(_6475_) );
	NAND2X1 NAND2X1_1313 ( .A(wSelec[138]), .B(_6475_), .Y(_6476_) );
	INVX1 INVX1_817 ( .A(wSelec[139]), .Y(_6477_) );
	NAND2X1 NAND2X1_1314 ( .A(wSelec[140]), .B(_6477_), .Y(_6478_) );
	NOR2X1 NOR2X1_753 ( .A(_6476_), .B(_6478_), .Y(_6479_) );
	NAND2X1 NAND2X1_1315 ( .A(wSelec[141]), .B(wSelec[142]), .Y(_6480_) );
	INVX1 INVX1_818 ( .A(_6480_), .Y(_6481_) );
	NAND2X1 NAND2X1_1316 ( .A(_6481_), .B(_6479_), .Y(_6482_) );
	INVX1 INVX1_819 ( .A(_6482_), .Y(_6483_) );
	AOI22X1 AOI22X1_1019 ( .A(_6474_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_6483_), .Y(_6484_) );
	OR2X2 OR2X2_74 ( .A(_6470_), .B(_6471_), .Y(_6485_) );
	OR2X2 OR2X2_75 ( .A(wSelec[141]), .B(wSelec[142]), .Y(_6486_) );
	NOR2X1 NOR2X1_754 ( .A(_6486_), .B(_6485_), .Y(_6487_) );
	NOR2X1 NOR2X1_755 ( .A(_6465_), .B(_6470_), .Y(_6488_) );
	INVX1 INVX1_820 ( .A(wSelec[141]), .Y(_6489_) );
	NAND2X1 NAND2X1_1317 ( .A(wSelec[142]), .B(_6489_), .Y(_6490_) );
	INVX2 INVX2_22 ( .A(_6490_), .Y(_6491_) );
	NAND2X1 NAND2X1_1318 ( .A(_6491_), .B(_6488_), .Y(_6492_) );
	INVX1 INVX1_821 ( .A(_6492_), .Y(_6493_) );
	AOI22X1 AOI22X1_1020 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_6487_), .C(_6493_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_6494_) );
	NAND3X1 NAND3X1_316 ( .A(_6468_), .B(_6494_), .C(_6484_), .Y(_6495_) );
	NOR2X1 NOR2X1_756 ( .A(wSelec[138]), .B(wSelec[137]), .Y(_6496_) );
	NOR2X1 NOR2X1_757 ( .A(wSelec[139]), .B(wSelec[140]), .Y(_6497_) );
	NAND2X1 NAND2X1_1319 ( .A(_6496_), .B(_6497_), .Y(_6498_) );
	NOR2X1 NOR2X1_758 ( .A(_6461_), .B(_6498_), .Y(_6499_) );
	NAND2X1 NAND2X1_1320 ( .A(wSelec[138]), .B(wSelec[137]), .Y(_6500_) );
	NOR3X1 NOR3X1_533 ( .A(_6471_), .B(_6500_), .C(_6461_), .Y(_6501_) );
	AOI22X1 AOI22X1_1021 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_6501_), .C(_6499_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_6502_) );
	INVX1 INVX1_822 ( .A(_6486_), .Y(_6503_) );
	NOR2X1 NOR2X1_759 ( .A(_6471_), .B(_6476_), .Y(_6504_) );
	AND2X2 AND2X2_143 ( .A(_6504_), .B(_6503_), .Y(_6505_) );
	NAND2X1 NAND2X1_1321 ( .A(wSelec[139]), .B(wSelec[140]), .Y(_6506_) );
	NOR3X1 NOR3X1_534 ( .A(_6480_), .B(_6500_), .C(_6506_), .Y(_6507_) );
	AOI22X1 AOI22X1_1022 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_6507_), .C(_6505_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_6508_) );
	INVX1 INVX1_823 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_6509_) );
	INVX1 INVX1_824 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_6510_) );
	NOR2X1 NOR2X1_760 ( .A(_6470_), .B(_6478_), .Y(_6511_) );
	NAND2X1 NAND2X1_1322 ( .A(_6481_), .B(_6511_), .Y(_6512_) );
	NOR2X1 NOR2X1_761 ( .A(_6500_), .B(_6506_), .Y(_6513_) );
	NAND2X1 NAND2X1_1323 ( .A(_6513_), .B(_6491_), .Y(_6514_) );
	OAI22X1 OAI22X1_173 ( .A(_6509_), .B(_6514_), .C(_6512_), .D(_6510_), .Y(_6515_) );
	INVX1 INVX1_825 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_6516_) );
	NOR3X1 NOR3X1_535 ( .A(_6461_), .B(_6476_), .C(_6478_), .Y(_6517_) );
	NAND2X1 NAND2X1_1324 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_6517_), .Y(_6518_) );
	NOR2X1 NOR2X1_762 ( .A(_6500_), .B(_6465_), .Y(_6519_) );
	NAND2X1 NAND2X1_1325 ( .A(_6491_), .B(_6519_), .Y(_6520_) );
	OAI21X1 OAI21X1_217 ( .A(_6516_), .B(_6520_), .C(_6518_), .Y(_6521_) );
	NOR2X1 NOR2X1_763 ( .A(_6515_), .B(_6521_), .Y(_6522_) );
	NAND3X1 NAND3X1_317 ( .A(_6502_), .B(_6508_), .C(_6522_), .Y(_6523_) );
	INVX1 INVX1_826 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_6524_) );
	INVX1 INVX1_827 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_6525_) );
	NOR2X1 NOR2X1_764 ( .A(_6465_), .B(_6476_), .Y(_6526_) );
	NAND2X1 NAND2X1_1326 ( .A(_6462_), .B(_6526_), .Y(_6527_) );
	NOR2X1 NOR2X1_765 ( .A(_6463_), .B(_6478_), .Y(_6528_) );
	NAND2X1 NAND2X1_1327 ( .A(_6462_), .B(_6528_), .Y(_6529_) );
	OAI22X1 OAI22X1_174 ( .A(_6529_), .B(_6524_), .C(_6525_), .D(_6527_), .Y(_6530_) );
	INVX1 INVX1_828 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_6531_) );
	INVX1 INVX1_829 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_6532_) );
	NAND2X1 NAND2X1_1328 ( .A(_6491_), .B(_6526_), .Y(_6533_) );
	NOR2X1 NOR2X1_766 ( .A(_6500_), .B(_6471_), .Y(_6534_) );
	NAND2X1 NAND2X1_1329 ( .A(_6491_), .B(_6534_), .Y(_6535_) );
	OAI22X1 OAI22X1_175 ( .A(_6531_), .B(_6535_), .C(_6533_), .D(_6532_), .Y(_6536_) );
	NOR2X1 NOR2X1_767 ( .A(_6536_), .B(_6530_), .Y(_6537_) );
	NOR3X1 NOR3X1_536 ( .A(_6470_), .B(_6506_), .C(_6490_), .Y(_6538_) );
	NAND2X1 NAND2X1_1330 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_6538_), .Y(_6539_) );
	NOR3X1 NOR3X1_537 ( .A(_6478_), .B(_6500_), .C(_6490_), .Y(_6540_) );
	NAND2X1 NAND2X1_1331 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_6540_), .Y(_6541_) );
	NAND2X1 NAND2X1_1332 ( .A(_6539_), .B(_6541_), .Y(_6542_) );
	INVX1 INVX1_830 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_6543_) );
	NAND2X1 NAND2X1_1333 ( .A(_6481_), .B(_6466_), .Y(_6544_) );
	NOR3X1 NOR3X1_538 ( .A(_6476_), .B(_6478_), .C(_6490_), .Y(_6545_) );
	NAND2X1 NAND2X1_1334 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_6545_), .Y(_6546_) );
	OAI21X1 OAI21X1_218 ( .A(_6543_), .B(_6544_), .C(_6546_), .Y(_6547_) );
	NOR2X1 NOR2X1_768 ( .A(_6542_), .B(_6547_), .Y(_6548_) );
	NAND2X1 NAND2X1_1335 ( .A(_6537_), .B(_6548_), .Y(_6549_) );
	NOR3X1 NOR3X1_539 ( .A(_6495_), .B(_6549_), .C(_6523_), .Y(_6550_) );
	NAND2X1 NAND2X1_1336 ( .A(_6462_), .B(_6519_), .Y(_6551_) );
	INVX1 INVX1_831 ( .A(_6551_), .Y(_6552_) );
	INVX1 INVX1_832 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_6553_) );
	NOR3X1 NOR3X1_540 ( .A(_6463_), .B(_6486_), .C(_6465_), .Y(_6554_) );
	NAND2X1 NAND2X1_1337 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_6554_), .Y(_6555_) );
	NAND2X1 NAND2X1_1338 ( .A(_6503_), .B(_6526_), .Y(_6556_) );
	OAI21X1 OAI21X1_219 ( .A(_6556_), .B(_6553_), .C(_6555_), .Y(_6557_) );
	AOI21X1 AOI21X1_155 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_6552_), .C(_6557_), .Y(_6558_) );
	INVX1 INVX1_833 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_6559_) );
	INVX1 INVX1_834 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_6560_) );
	NOR2X1 NOR2X1_769 ( .A(_6506_), .B(_6463_), .Y(_6561_) );
	NAND2X1 NAND2X1_1339 ( .A(_6462_), .B(_6561_), .Y(_6562_) );
	NAND2X1 NAND2X1_1340 ( .A(_6503_), .B(_6488_), .Y(_6563_) );
	OAI22X1 OAI22X1_176 ( .A(_6560_), .B(_6562_), .C(_6563_), .D(_6559_), .Y(_6564_) );
	INVX1 INVX1_835 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_6565_) );
	INVX1 INVX1_836 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_6566_) );
	NAND2X1 NAND2X1_1341 ( .A(_6462_), .B(_6488_), .Y(_6567_) );
	NAND2X1 NAND2X1_1342 ( .A(_6503_), .B(_6534_), .Y(_6568_) );
	OAI22X1 OAI22X1_177 ( .A(_6565_), .B(_6568_), .C(_6567_), .D(_6566_), .Y(_6569_) );
	NOR2X1 NOR2X1_770 ( .A(_6564_), .B(_6569_), .Y(_6570_) );
	INVX1 INVX1_837 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_6571_) );
	NOR3X1 NOR3X1_541 ( .A(_6486_), .B(_6500_), .C(_6465_), .Y(_6572_) );
	NAND2X1 NAND2X1_1343 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_6572_), .Y(_6573_) );
	OR2X2 OR2X2_76 ( .A(_6498_), .B(_6480_), .Y(_6574_) );
	OAI21X1 OAI21X1_220 ( .A(_6571_), .B(_6574_), .C(_6573_), .Y(_6575_) );
	INVX1 INVX1_838 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_6576_) );
	INVX1 INVX1_839 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_6577_) );
	NOR2X1 NOR2X1_771 ( .A(_6506_), .B(_6476_), .Y(_6578_) );
	NAND2X1 NAND2X1_1344 ( .A(_6462_), .B(_6578_), .Y(_6579_) );
	NAND2X1 NAND2X1_1345 ( .A(_6481_), .B(_6472_), .Y(_6580_) );
	OAI22X1 OAI22X1_178 ( .A(_6579_), .B(_6577_), .C(_6576_), .D(_6580_), .Y(_6581_) );
	NOR2X1 NOR2X1_772 ( .A(_6575_), .B(_6581_), .Y(_6582_) );
	NAND3X1 NAND3X1_318 ( .A(_6558_), .B(_6582_), .C(_6570_), .Y(_6583_) );
	NOR3X1 NOR3X1_542 ( .A(_6463_), .B(_6471_), .C(_6486_), .Y(_6584_) );
	NOR3X1 NOR3X1_543 ( .A(_6480_), .B(_6506_), .C(_6470_), .Y(_6585_) );
	AOI22X1 AOI22X1_1023 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_6584_), .C(_6585_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_6586_) );
	NOR3X1 NOR3X1_544 ( .A(_6480_), .B(_6506_), .C(_6476_), .Y(_6587_) );
	NOR3X1 NOR3X1_545 ( .A(_6480_), .B(_6500_), .C(_6478_), .Y(_6588_) );
	AOI22X1 AOI22X1_1024 ( .A(_6587_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_6588_), .Y(_6589_) );
	NAND2X1 NAND2X1_1346 ( .A(_6586_), .B(_6589_), .Y(_6590_) );
	NOR3X1 NOR3X1_546 ( .A(_6478_), .B(_6463_), .C(_6490_), .Y(_6591_) );
	NOR3X1 NOR3X1_547 ( .A(_6470_), .B(_6478_), .C(_6490_), .Y(_6592_) );
	AOI22X1 AOI22X1_1025 ( .A(_6591_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_6592_), .Y(_6593_) );
	NOR3X1 NOR3X1_548 ( .A(_6461_), .B(_6506_), .C(_6470_), .Y(_6594_) );
	NOR3X1 NOR3X1_549 ( .A(_6500_), .B(_6506_), .C(_6461_), .Y(_6595_) );
	AOI22X1 AOI22X1_1026 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_6595_), .C(_6594_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_6596_) );
	NAND2X1 NAND2X1_1347 ( .A(_6596_), .B(_6593_), .Y(_6597_) );
	NOR2X1 NOR2X1_773 ( .A(_6590_), .B(_6597_), .Y(_6598_) );
	NOR3X1 NOR3X1_550 ( .A(_6486_), .B(_6506_), .C(_6470_), .Y(_6599_) );
	NOR3X1 NOR3X1_551 ( .A(_6486_), .B(_6506_), .C(_6476_), .Y(_6600_) );
	AOI22X1 AOI22X1_1027 ( .A(_6599_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_6600_), .Y(_6601_) );
	NOR3X1 NOR3X1_552 ( .A(_6486_), .B(_6500_), .C(_6478_), .Y(_6602_) );
	NOR3X1 NOR3X1_553 ( .A(_6461_), .B(_6471_), .C(_6476_), .Y(_6603_) );
	AOI22X1 AOI22X1_1028 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_6602_), .C(_6603_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_6604_) );
	NAND2X1 NAND2X1_1348 ( .A(_6601_), .B(_6604_), .Y(_6605_) );
	NOR3X1 NOR3X1_554 ( .A(_6500_), .B(_6506_), .C(_6486_), .Y(_6606_) );
	NOR3X1 NOR3X1_555 ( .A(_6476_), .B(_6471_), .C(_6490_), .Y(_6607_) );
	AOI22X1 AOI22X1_1029 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_6606_), .C(_6607_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_6608_) );
	NOR3X1 NOR3X1_556 ( .A(_6463_), .B(_6471_), .C(_6490_), .Y(_6609_) );
	NOR3X1 NOR3X1_557 ( .A(_6463_), .B(_6506_), .C(_6490_), .Y(_6610_) );
	AOI22X1 AOI22X1_1030 ( .A(_6609_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_6610_), .Y(_6611_) );
	NAND2X1 NAND2X1_1349 ( .A(_6611_), .B(_6608_), .Y(_6612_) );
	NOR2X1 NOR2X1_774 ( .A(_6605_), .B(_6612_), .Y(_6613_) );
	NAND2X1 NAND2X1_1350 ( .A(_6613_), .B(_6598_), .Y(_6614_) );
	NOR3X1 NOR3X1_558 ( .A(_6461_), .B(_6500_), .C(_6478_), .Y(_6615_) );
	NOR3X1 NOR3X1_559 ( .A(_6471_), .B(_6480_), .C(_6476_), .Y(_6616_) );
	AOI22X1 AOI22X1_1031 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_6616_), .C(_6615_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_6617_) );
	NOR3X1 NOR3X1_560 ( .A(_6465_), .B(_6463_), .C(_6490_), .Y(_6618_) );
	NOR3X1 NOR3X1_561 ( .A(_6476_), .B(_6506_), .C(_6490_), .Y(_6619_) );
	AOI22X1 AOI22X1_1032 ( .A(_6618_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_6619_), .Y(_6620_) );
	NAND2X1 NAND2X1_1351 ( .A(_6617_), .B(_6620_), .Y(_6621_) );
	NOR3X1 NOR3X1_562 ( .A(_6461_), .B(_6470_), .C(_6478_), .Y(_6622_) );
	NAND2X1 NAND2X1_1352 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_6622_), .Y(_6623_) );
	NOR3X1 NOR3X1_563 ( .A(_6480_), .B(_6500_), .C(_6465_), .Y(_6624_) );
	NAND2X1 NAND2X1_1353 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_6624_), .Y(_6625_) );
	NOR3X1 NOR3X1_564 ( .A(_6463_), .B(_6506_), .C(_6486_), .Y(_6626_) );
	NOR3X1 NOR3X1_565 ( .A(_6463_), .B(_6480_), .C(_6478_), .Y(_6627_) );
	AOI22X1 AOI22X1_1033 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_6626_), .C(_6627_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_6628_) );
	NAND3X1 NAND3X1_319 ( .A(_6623_), .B(_6625_), .C(_6628_), .Y(_6629_) );
	NOR2X1 NOR2X1_775 ( .A(_6629_), .B(_6621_), .Y(_6630_) );
	NOR3X1 NOR3X1_566 ( .A(_6463_), .B(_6486_), .C(_6478_), .Y(_6631_) );
	NOR3X1 NOR3X1_567 ( .A(_6465_), .B(_6480_), .C(_6470_), .Y(_6632_) );
	AOI22X1 AOI22X1_1034 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_6631_), .C(_6632_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_6633_) );
	NOR3X1 NOR3X1_568 ( .A(_6465_), .B(_6480_), .C(_6476_), .Y(_6634_) );
	NAND2X1 NAND2X1_1354 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_6634_), .Y(_6635_) );
	NOR3X1 NOR3X1_569 ( .A(_6470_), .B(_6471_), .C(_6490_), .Y(_6636_) );
	NAND2X1 NAND2X1_1355 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_6636_), .Y(_6637_) );
	NAND3X1 NAND3X1_320 ( .A(_6635_), .B(_6637_), .C(_6633_), .Y(_6638_) );
	NOR3X1 NOR3X1_570 ( .A(_6470_), .B(_6486_), .C(_6478_), .Y(_6639_) );
	NOR3X1 NOR3X1_571 ( .A(_6480_), .B(_6506_), .C(_6463_), .Y(_6640_) );
	AOI22X1 AOI22X1_1035 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_6640_), .C(_6639_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_6641_) );
	NOR3X1 NOR3X1_572 ( .A(_6476_), .B(_6486_), .C(_6478_), .Y(_6642_) );
	NOR3X1 NOR3X1_573 ( .A(_6480_), .B(_6500_), .C(_6471_), .Y(_6643_) );
	AOI22X1 AOI22X1_1036 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_6643_), .C(_6642_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_6644_) );
	NAND2X1 NAND2X1_1356 ( .A(_6641_), .B(_6644_), .Y(_6645_) );
	NOR2X1 NOR2X1_776 ( .A(_6645_), .B(_6638_), .Y(_6646_) );
	NAND2X1 NAND2X1_1357 ( .A(_6630_), .B(_6646_), .Y(_6647_) );
	NOR3X1 NOR3X1_574 ( .A(_6614_), .B(_6583_), .C(_6647_), .Y(_6648_) );
	INVX1 INVX1_840 ( .A(wSelec[134]), .Y(_6649_) );
	NAND2X1 NAND2X1_1358 ( .A(wSelec[133]), .B(_6649_), .Y(_6650_) );
	INVX1 INVX1_841 ( .A(wSelec[136]), .Y(_6651_) );
	NAND2X1 NAND2X1_1359 ( .A(wSelec[135]), .B(_6651_), .Y(_6652_) );
	NOR2X1 NOR2X1_777 ( .A(_6650_), .B(_6652_), .Y(_6653_) );
	NOR2X1 NOR2X1_778 ( .A(wSelec[134]), .B(wSelec[133]), .Y(_6654_) );
	INVX1 INVX1_842 ( .A(_6654_), .Y(_6655_) );
	NOR2X1 NOR2X1_779 ( .A(_6652_), .B(_6655_), .Y(_6656_) );
	AOI22X1 AOI22X1_1037 ( .A(wData[20]), .B(_6653_), .C(_6656_), .D(wData[16]), .Y(_6657_) );
	INVX1 INVX1_843 ( .A(wSelec[133]), .Y(_6658_) );
	NAND2X1 NAND2X1_1360 ( .A(wSelec[134]), .B(_6658_), .Y(_6659_) );
	NOR2X1 NOR2X1_780 ( .A(_6659_), .B(_6652_), .Y(_6660_) );
	NAND2X1 NAND2X1_1361 ( .A(wData[24]), .B(_6660_), .Y(_6661_) );
	INVX1 INVX1_844 ( .A(wSelec[135]), .Y(_6662_) );
	NAND2X1 NAND2X1_1362 ( .A(_6662_), .B(_6651_), .Y(_6663_) );
	NOR2X1 NOR2X1_781 ( .A(_6650_), .B(_6663_), .Y(_6664_) );
	NAND2X1 NAND2X1_1363 ( .A(wSelec[134]), .B(wSelec[133]), .Y(_6665_) );
	NOR2X1 NOR2X1_782 ( .A(_6665_), .B(_6652_), .Y(_6666_) );
	AOI22X1 AOI22X1_1038 ( .A(_6666_), .B(wData[28]), .C(wData[4]), .D(_6664_), .Y(_6667_) );
	NAND3X1 NAND3X1_321 ( .A(_6661_), .B(_6667_), .C(_6657_), .Y(_6668_) );
	NAND2X1 NAND2X1_1364 ( .A(wSelec[136]), .B(_6662_), .Y(_6669_) );
	NOR2X1 NOR2X1_783 ( .A(_6669_), .B(_6655_), .Y(_6670_) );
	NAND2X1 NAND2X1_1365 ( .A(wData[32]), .B(_6670_), .Y(_6671_) );
	NAND2X1 NAND2X1_1366 ( .A(wSelec[135]), .B(wSelec[136]), .Y(_6672_) );
	NOR2X1 NOR2X1_784 ( .A(_6672_), .B(_6659_), .Y(_6673_) );
	NOR2X1 NOR2X1_785 ( .A(_6672_), .B(_6650_), .Y(_6674_) );
	AOI22X1 AOI22X1_1039 ( .A(_6673_), .B(wData[56]), .C(wData[52]), .D(_6674_), .Y(_6675_) );
	NOR2X1 NOR2X1_786 ( .A(_6665_), .B(_6672_), .Y(_6676_) );
	NOR2X1 NOR2X1_787 ( .A(_6665_), .B(_6669_), .Y(_6677_) );
	AOI22X1 AOI22X1_1040 ( .A(wData[60]), .B(_6676_), .C(_6677_), .D(wData[44]), .Y(_6678_) );
	NAND3X1 NAND3X1_322 ( .A(_6671_), .B(_6678_), .C(_6675_), .Y(_6679_) );
	NOR2X1 NOR2X1_788 ( .A(_6659_), .B(_6669_), .Y(_6680_) );
	NAND2X1 NAND2X1_1367 ( .A(wData[40]), .B(_6680_), .Y(_6681_) );
	NOR2X1 NOR2X1_789 ( .A(_6669_), .B(_6650_), .Y(_6682_) );
	NAND2X1 NAND2X1_1368 ( .A(wData[36]), .B(_6682_), .Y(_6683_) );
	NOR2X1 NOR2X1_790 ( .A(_6663_), .B(_6655_), .Y(_6684_) );
	NAND2X1 NAND2X1_1369 ( .A(wData[0]), .B(_6684_), .Y(_6685_) );
	NAND3X1 NAND3X1_323 ( .A(_6681_), .B(_6683_), .C(_6685_), .Y(_6686_) );
	INVX1 INVX1_845 ( .A(wData[48]), .Y(_6687_) );
	NOR2X1 NOR2X1_791 ( .A(_6662_), .B(_6651_), .Y(_6688_) );
	NAND2X1 NAND2X1_1370 ( .A(_6654_), .B(_6688_), .Y(_6689_) );
	NOR2X1 NOR2X1_792 ( .A(_6659_), .B(_6663_), .Y(_6690_) );
	NOR2X1 NOR2X1_793 ( .A(_6665_), .B(_6663_), .Y(_6691_) );
	AOI22X1 AOI22X1_1041 ( .A(_6690_), .B(wData[8]), .C(wData[12]), .D(_6691_), .Y(_6692_) );
	OAI21X1 OAI21X1_221 ( .A(_6687_), .B(_6689_), .C(_6692_), .Y(_6693_) );
	OR2X2 OR2X2_77 ( .A(_6693_), .B(_6686_), .Y(_6694_) );
	NOR3X1 NOR3X1_575 ( .A(_6668_), .B(_6679_), .C(_6694_), .Y(_6695_) );
	AND2X2 AND2X2_144 ( .A(_6695_), .B(_6459_), .Y(_6696_) );
	AOI21X1 AOI21X1_156 ( .A(_6550_), .B(_6648_), .C(_6696_), .Y(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_0_) );
	INVX1 INVX1_846 ( .A(_6567_), .Y(_6697_) );
	AOI21X1 AOI21X1_157 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_6697_), .C(_6459_), .Y(_6698_) );
	AOI22X1 AOI22X1_1042 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_6467_), .C(_6483_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_6699_) );
	AOI22X1 AOI22X1_1043 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_6487_), .C(_6493_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_6700_) );
	NAND3X1 NAND3X1_324 ( .A(_6698_), .B(_6699_), .C(_6700_), .Y(_6701_) );
	INVX1 INVX1_847 ( .A(_6527_), .Y(_6702_) );
	AOI22X1 AOI22X1_1044 ( .A(_6552_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_6702_), .Y(_6703_) );
	AOI22X1 AOI22X1_1045 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_6626_), .C(_6505_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_6704_) );
	INVX1 INVX1_848 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_6705_) );
	INVX1 INVX1_849 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_6706_) );
	OAI22X1 OAI22X1_179 ( .A(_6705_), .B(_6514_), .C(_6512_), .D(_6706_), .Y(_6707_) );
	INVX1 INVX1_850 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_6708_) );
	NAND2X1 NAND2X1_1371 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_6615_), .Y(_6709_) );
	OAI21X1 OAI21X1_222 ( .A(_6708_), .B(_6520_), .C(_6709_), .Y(_6710_) );
	NOR2X1 NOR2X1_794 ( .A(_6707_), .B(_6710_), .Y(_6711_) );
	NAND3X1 NAND3X1_325 ( .A(_6703_), .B(_6704_), .C(_6711_), .Y(_6712_) );
	INVX1 INVX1_851 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_6713_) );
	NAND2X1 NAND2X1_1372 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_6499_), .Y(_6714_) );
	OAI21X1 OAI21X1_223 ( .A(_6713_), .B(_6529_), .C(_6714_), .Y(_6715_) );
	INVX1 INVX1_852 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_6716_) );
	INVX1 INVX1_853 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_6717_) );
	OAI22X1 OAI22X1_180 ( .A(_6716_), .B(_6535_), .C(_6533_), .D(_6717_), .Y(_6718_) );
	NOR2X1 NOR2X1_795 ( .A(_6718_), .B(_6715_), .Y(_6719_) );
	AOI22X1 AOI22X1_1046 ( .A(_6619_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_6592_), .Y(_6720_) );
	AND2X2 AND2X2_145 ( .A(_6466_), .B(_6481_), .Y(_6721_) );
	AOI22X1 AOI22X1_1047 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_6591_), .C(_6721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_6722_) );
	NAND3X1 NAND3X1_326 ( .A(_6720_), .B(_6722_), .C(_6719_), .Y(_6723_) );
	NOR3X1 NOR3X1_576 ( .A(_6723_), .B(_6701_), .C(_6712_), .Y(_6724_) );
	INVX1 INVX1_854 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_6725_) );
	NAND2X1 NAND2X1_1373 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_6554_), .Y(_6726_) );
	OAI21X1 OAI21X1_224 ( .A(_6556_), .B(_6725_), .C(_6726_), .Y(_6727_) );
	AOI21X1 AOI21X1_158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_6603_), .C(_6727_), .Y(_6728_) );
	INVX1 INVX1_855 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_6729_) );
	INVX1 INVX1_856 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_6730_) );
	OAI22X1 OAI22X1_181 ( .A(_6730_), .B(_6562_), .C(_6563_), .D(_6729_), .Y(_6731_) );
	INVX1 INVX1_857 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_6732_) );
	NAND2X1 NAND2X1_1374 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_6572_), .Y(_6733_) );
	OAI21X1 OAI21X1_225 ( .A(_6473_), .B(_6732_), .C(_6733_), .Y(_6734_) );
	NOR2X1 NOR2X1_796 ( .A(_6734_), .B(_6731_), .Y(_6735_) );
	INVX1 INVX1_858 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_6736_) );
	INVX1 INVX1_859 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_6737_) );
	OAI22X1 OAI22X1_182 ( .A(_6568_), .B(_6737_), .C(_6574_), .D(_6736_), .Y(_6738_) );
	INVX1 INVX1_860 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_6739_) );
	NOR2X1 NOR2X1_797 ( .A(_6739_), .B(_6579_), .Y(_6740_) );
	INVX1 INVX1_861 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_6741_) );
	NOR2X1 NOR2X1_798 ( .A(_6741_), .B(_6580_), .Y(_6742_) );
	NOR3X1 NOR3X1_577 ( .A(_6740_), .B(_6738_), .C(_6742_), .Y(_6743_) );
	NAND3X1 NAND3X1_327 ( .A(_6735_), .B(_6728_), .C(_6743_), .Y(_6744_) );
	AOI22X1 AOI22X1_1048 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_6584_), .C(_6585_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_6745_) );
	AOI22X1 AOI22X1_1049 ( .A(_6587_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_6588_), .Y(_6746_) );
	NAND2X1 NAND2X1_1375 ( .A(_6745_), .B(_6746_), .Y(_6747_) );
	AOI22X1 AOI22X1_1050 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_6595_), .C(_6594_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_6748_) );
	AOI22X1 AOI22X1_1051 ( .A(_6538_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_6545_), .Y(_6749_) );
	NAND2X1 NAND2X1_1376 ( .A(_6748_), .B(_6749_), .Y(_6750_) );
	NOR2X1 NOR2X1_799 ( .A(_6747_), .B(_6750_), .Y(_6751_) );
	AOI22X1 AOI22X1_1052 ( .A(_6599_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_6600_), .Y(_6752_) );
	AOI22X1 AOI22X1_1053 ( .A(_6501_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_6602_), .Y(_6753_) );
	NAND2X1 NAND2X1_1377 ( .A(_6752_), .B(_6753_), .Y(_6754_) );
	AOI22X1 AOI22X1_1054 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_6606_), .C(_6607_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_6755_) );
	AOI22X1 AOI22X1_1055 ( .A(_6609_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_6610_), .Y(_6756_) );
	NAND2X1 NAND2X1_1378 ( .A(_6756_), .B(_6755_), .Y(_6757_) );
	NOR2X1 NOR2X1_800 ( .A(_6754_), .B(_6757_), .Y(_6758_) );
	NAND2X1 NAND2X1_1379 ( .A(_6758_), .B(_6751_), .Y(_6759_) );
	AOI22X1 AOI22X1_1056 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_6616_), .C(_6517_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_6760_) );
	AOI22X1 AOI22X1_1057 ( .A(_6540_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_6618_), .Y(_6761_) );
	NAND2X1 NAND2X1_1380 ( .A(_6760_), .B(_6761_), .Y(_6762_) );
	AOI22X1 AOI22X1_1058 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_6507_), .C(_6627_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_6763_) );
	NAND2X1 NAND2X1_1381 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_6622_), .Y(_6764_) );
	NAND2X1 NAND2X1_1382 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_6624_), .Y(_6765_) );
	NAND3X1 NAND3X1_328 ( .A(_6764_), .B(_6765_), .C(_6763_), .Y(_6766_) );
	NOR2X1 NOR2X1_801 ( .A(_6766_), .B(_6762_), .Y(_6767_) );
	AOI22X1 AOI22X1_1059 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_6631_), .C(_6632_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_6768_) );
	NAND2X1 NAND2X1_1383 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_6634_), .Y(_6769_) );
	NAND2X1 NAND2X1_1384 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_6636_), .Y(_6770_) );
	NAND3X1 NAND3X1_329 ( .A(_6769_), .B(_6770_), .C(_6768_), .Y(_6771_) );
	AOI22X1 AOI22X1_1060 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_6640_), .C(_6639_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_6772_) );
	AOI22X1 AOI22X1_1061 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_6643_), .C(_6642_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_6773_) );
	NAND2X1 NAND2X1_1385 ( .A(_6772_), .B(_6773_), .Y(_6774_) );
	NOR2X1 NOR2X1_802 ( .A(_6774_), .B(_6771_), .Y(_6775_) );
	NAND2X1 NAND2X1_1386 ( .A(_6767_), .B(_6775_), .Y(_6776_) );
	NOR3X1 NOR3X1_578 ( .A(_6759_), .B(_6744_), .C(_6776_), .Y(_6777_) );
	AOI21X1 AOI21X1_159 ( .A(wData[21]), .B(_6653_), .C(_6458_), .Y(_6778_) );
	AOI22X1 AOI22X1_1062 ( .A(_6656_), .B(wData[17]), .C(wData[1]), .D(_6684_), .Y(_6779_) );
	AOI22X1 AOI22X1_1063 ( .A(_6677_), .B(wData[45]), .C(wData[25]), .D(_6660_), .Y(_6780_) );
	NAND3X1 NAND3X1_330 ( .A(_6778_), .B(_6780_), .C(_6779_), .Y(_6781_) );
	NAND3X1 NAND3X1_331 ( .A(wData[49]), .B(_6654_), .C(_6688_), .Y(_6782_) );
	AOI22X1 AOI22X1_1064 ( .A(wData[61]), .B(_6676_), .C(_6664_), .D(wData[5]), .Y(_6783_) );
	AND2X2 AND2X2_146 ( .A(_6783_), .B(_6782_), .Y(_6784_) );
	AOI22X1 AOI22X1_1065 ( .A(_6673_), .B(wData[57]), .C(wData[41]), .D(_6680_), .Y(_6785_) );
	AOI22X1 AOI22X1_1066 ( .A(wData[53]), .B(_6674_), .C(_6670_), .D(wData[33]), .Y(_6786_) );
	AND2X2 AND2X2_147 ( .A(_6786_), .B(_6785_), .Y(_6787_) );
	AOI22X1 AOI22X1_1067 ( .A(_6690_), .B(wData[9]), .C(wData[13]), .D(_6691_), .Y(_6788_) );
	AOI22X1 AOI22X1_1068 ( .A(_6666_), .B(wData[29]), .C(wData[37]), .D(_6682_), .Y(_6789_) );
	AND2X2 AND2X2_148 ( .A(_6788_), .B(_6789_), .Y(_6790_) );
	NAND3X1 NAND3X1_332 ( .A(_6784_), .B(_6790_), .C(_6787_), .Y(_6791_) );
	NOR2X1 NOR2X1_803 ( .A(_6781_), .B(_6791_), .Y(_6792_) );
	AOI21X1 AOI21X1_160 ( .A(_6724_), .B(_6777_), .C(_6792_), .Y(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_1_) );
	AOI21X1 AOI21X1_161 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_6697_), .C(_6459_), .Y(_6793_) );
	INVX1 INVX1_862 ( .A(_6556_), .Y(_6794_) );
	AOI22X1 AOI22X1_1069 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_6467_), .C(_6794_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_6795_) );
	INVX1 INVX1_863 ( .A(_6568_), .Y(_6796_) );
	AOI22X1 AOI22X1_1070 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_6603_), .C(_6796_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_6797_) );
	NAND3X1 NAND3X1_333 ( .A(_6797_), .B(_6793_), .C(_6795_), .Y(_6798_) );
	AOI22X1 AOI22X1_1071 ( .A(_6552_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_6702_), .Y(_6799_) );
	AOI22X1 AOI22X1_1072 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_6501_), .C(_6474_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_6800_) );
	INVX1 INVX1_864 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_6801_) );
	NAND2X1 NAND2X1_1387 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_6591_), .Y(_6802_) );
	OAI21X1 OAI21X1_226 ( .A(_6801_), .B(_6563_), .C(_6802_), .Y(_6803_) );
	INVX1 INVX1_865 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_6804_) );
	NAND2X1 NAND2X1_1388 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_6517_), .Y(_6805_) );
	OAI21X1 OAI21X1_227 ( .A(_6804_), .B(_6520_), .C(_6805_), .Y(_6806_) );
	NOR2X1 NOR2X1_804 ( .A(_6803_), .B(_6806_), .Y(_6807_) );
	NAND3X1 NAND3X1_334 ( .A(_6799_), .B(_6800_), .C(_6807_), .Y(_6808_) );
	INVX1 INVX1_866 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_6809_) );
	NAND2X1 NAND2X1_1389 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_6499_), .Y(_6810_) );
	OAI21X1 OAI21X1_228 ( .A(_6809_), .B(_6529_), .C(_6810_), .Y(_6811_) );
	INVX1 INVX1_867 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_6812_) );
	INVX1 INVX1_868 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_6813_) );
	OAI22X1 OAI22X1_183 ( .A(_6812_), .B(_6535_), .C(_6533_), .D(_6813_), .Y(_6814_) );
	NOR2X1 NOR2X1_805 ( .A(_6814_), .B(_6811_), .Y(_6815_) );
	AOI22X1 AOI22X1_1073 ( .A(_6619_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_6592_), .Y(_6816_) );
	AND2X2 AND2X2_149 ( .A(_6491_), .B(_6513_), .Y(_6817_) );
	AOI22X1 AOI22X1_1074 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_6817_), .C(_6721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_6818_) );
	NAND3X1 NAND3X1_335 ( .A(_6816_), .B(_6818_), .C(_6815_), .Y(_6819_) );
	NOR3X1 NOR3X1_579 ( .A(_6819_), .B(_6798_), .C(_6808_), .Y(_6820_) );
	INVX1 INVX1_869 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_6821_) );
	NOR3X1 NOR3X1_580 ( .A(_6821_), .B(_6486_), .C(_6485_), .Y(_6822_) );
	AND2X2 AND2X2_150 ( .A(_6507_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_6823_) );
	AND2X2 AND2X2_151 ( .A(_6627_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_6824_) );
	NOR3X1 NOR3X1_581 ( .A(_6824_), .B(_6823_), .C(_6822_), .Y(_6825_) );
	INVX1 INVX1_870 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_6826_) );
	INVX1 INVX1_871 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_6827_) );
	OAI22X1 OAI22X1_184 ( .A(_6827_), .B(_6562_), .C(_6512_), .D(_6826_), .Y(_6828_) );
	INVX1 INVX1_872 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_6829_) );
	INVX1 INVX1_873 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_6830_) );
	NAND2X1 NAND2X1_1390 ( .A(_6503_), .B(_6504_), .Y(_6831_) );
	OAI22X1 OAI22X1_185 ( .A(_6831_), .B(_6830_), .C(_6829_), .D(_6482_), .Y(_6832_) );
	NOR2X1 NOR2X1_806 ( .A(_6828_), .B(_6832_), .Y(_6833_) );
	INVX1 INVX1_874 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_6834_) );
	NOR3X1 NOR3X1_582 ( .A(_6463_), .B(_6480_), .C(_6471_), .Y(_6835_) );
	NAND2X1 NAND2X1_1391 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_6835_), .Y(_6836_) );
	OAI21X1 OAI21X1_229 ( .A(_6492_), .B(_6834_), .C(_6836_), .Y(_6837_) );
	INVX1 INVX1_875 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_6838_) );
	INVX1 INVX1_876 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_6839_) );
	OAI22X1 OAI22X1_186 ( .A(_6579_), .B(_6839_), .C(_6838_), .D(_6580_), .Y(_6840_) );
	NOR2X1 NOR2X1_807 ( .A(_6837_), .B(_6840_), .Y(_6841_) );
	NAND3X1 NAND3X1_336 ( .A(_6825_), .B(_6841_), .C(_6833_), .Y(_6842_) );
	AOI22X1 AOI22X1_1075 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_6584_), .C(_6585_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_6843_) );
	AOI22X1 AOI22X1_1076 ( .A(_6587_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_6588_), .Y(_6844_) );
	NAND2X1 NAND2X1_1392 ( .A(_6843_), .B(_6844_), .Y(_6845_) );
	AOI22X1 AOI22X1_1077 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_6595_), .C(_6594_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_6846_) );
	AOI22X1 AOI22X1_1078 ( .A(_6538_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_6545_), .Y(_6847_) );
	NAND2X1 NAND2X1_1393 ( .A(_6846_), .B(_6847_), .Y(_6848_) );
	NOR2X1 NOR2X1_808 ( .A(_6845_), .B(_6848_), .Y(_6849_) );
	AOI22X1 AOI22X1_1079 ( .A(_6599_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_6600_), .Y(_6850_) );
	AOI22X1 AOI22X1_1080 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_6626_), .C(_6602_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_6851_) );
	NAND2X1 NAND2X1_1394 ( .A(_6851_), .B(_6850_), .Y(_6852_) );
	AOI22X1 AOI22X1_1081 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_6606_), .C(_6607_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_6853_) );
	AOI22X1 AOI22X1_1082 ( .A(_6609_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_6610_), .Y(_6854_) );
	NAND2X1 NAND2X1_1395 ( .A(_6854_), .B(_6853_), .Y(_6855_) );
	NOR2X1 NOR2X1_809 ( .A(_6852_), .B(_6855_), .Y(_6856_) );
	NAND2X1 NAND2X1_1396 ( .A(_6856_), .B(_6849_), .Y(_6857_) );
	AOI22X1 AOI22X1_1083 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_6616_), .C(_6615_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_6858_) );
	AOI22X1 AOI22X1_1084 ( .A(_6540_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_6618_), .Y(_6859_) );
	NAND2X1 NAND2X1_1397 ( .A(_6858_), .B(_6859_), .Y(_6860_) );
	AOI22X1 AOI22X1_1085 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_6624_), .C(_6622_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_6861_) );
	AOI22X1 AOI22X1_1086 ( .A(_6554_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_6572_), .Y(_6862_) );
	NAND2X1 NAND2X1_1398 ( .A(_6862_), .B(_6861_), .Y(_6863_) );
	NOR2X1 NOR2X1_810 ( .A(_6863_), .B(_6860_), .Y(_6864_) );
	AOI22X1 AOI22X1_1087 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_6631_), .C(_6632_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_6865_) );
	NAND2X1 NAND2X1_1399 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_6634_), .Y(_6866_) );
	NAND2X1 NAND2X1_1400 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_6636_), .Y(_6867_) );
	NAND3X1 NAND3X1_337 ( .A(_6866_), .B(_6867_), .C(_6865_), .Y(_6868_) );
	AOI22X1 AOI22X1_1088 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_6640_), .C(_6639_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_6869_) );
	AOI22X1 AOI22X1_1089 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_6643_), .C(_6642_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_6870_) );
	NAND2X1 NAND2X1_1401 ( .A(_6869_), .B(_6870_), .Y(_6871_) );
	NOR2X1 NOR2X1_811 ( .A(_6871_), .B(_6868_), .Y(_6872_) );
	NAND2X1 NAND2X1_1402 ( .A(_6864_), .B(_6872_), .Y(_6873_) );
	NOR3X1 NOR3X1_583 ( .A(_6857_), .B(_6842_), .C(_6873_), .Y(_6874_) );
	AOI22X1 AOI22X1_1090 ( .A(_6680_), .B(wData[42]), .C(wData[38]), .D(_6682_), .Y(_6875_) );
	AOI22X1 AOI22X1_1091 ( .A(_6677_), .B(wData[46]), .C(_6684_), .D(wData[2]), .Y(_6876_) );
	NAND2X1 NAND2X1_1403 ( .A(_6875_), .B(_6876_), .Y(_6877_) );
	AOI21X1 AOI21X1_162 ( .A(wData[34]), .B(_6670_), .C(_6877_), .Y(_6878_) );
	INVX1 INVX1_877 ( .A(wData[50]), .Y(_6879_) );
	AOI22X1 AOI22X1_1092 ( .A(_6690_), .B(wData[10]), .C(wData[14]), .D(_6691_), .Y(_6880_) );
	OAI21X1 OAI21X1_230 ( .A(_6879_), .B(_6689_), .C(_6880_), .Y(_6881_) );
	AOI22X1 AOI22X1_1093 ( .A(_6653_), .B(wData[22]), .C(wData[18]), .D(_6656_), .Y(_6882_) );
	NAND2X1 NAND2X1_1404 ( .A(wData[26]), .B(_6660_), .Y(_6883_) );
	AOI22X1 AOI22X1_1094 ( .A(_6666_), .B(wData[30]), .C(wData[6]), .D(_6664_), .Y(_6884_) );
	NAND3X1 NAND3X1_338 ( .A(_6883_), .B(_6884_), .C(_6882_), .Y(_6885_) );
	NOR2X1 NOR2X1_812 ( .A(_6881_), .B(_6885_), .Y(_6886_) );
	NAND2X1 NAND2X1_1405 ( .A(wData[58]), .B(_6673_), .Y(_6887_) );
	NAND2X1 NAND2X1_1406 ( .A(wData[54]), .B(_6674_), .Y(_6888_) );
	NAND2X1 NAND2X1_1407 ( .A(_6887_), .B(_6888_), .Y(_6889_) );
	AOI21X1 AOI21X1_163 ( .A(wData[62]), .B(_6676_), .C(_6889_), .Y(_6890_) );
	NAND3X1 NAND3X1_339 ( .A(_6878_), .B(_6890_), .C(_6886_), .Y(_6891_) );
	NOR2X1 NOR2X1_813 ( .A(_6458_), .B(_6891_), .Y(_6892_) );
	AOI21X1 AOI21X1_164 ( .A(_6820_), .B(_6874_), .C(_6892_), .Y(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_2_) );
	AOI21X1 AOI21X1_165 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_6702_), .C(_6459_), .Y(_6893_) );
	AOI22X1 AOI22X1_1095 ( .A(_6474_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_6794_), .Y(_6894_) );
	AOI22X1 AOI22X1_1096 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_6796_), .C(_6552_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_6895_) );
	NAND3X1 NAND3X1_340 ( .A(_6895_), .B(_6893_), .C(_6894_), .Y(_6896_) );
	AOI22X1 AOI22X1_1097 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_6501_), .C(_6499_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_6897_) );
	AOI22X1 AOI22X1_1098 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_6572_), .C(_6697_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_6898_) );
	INVX1 INVX1_878 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_6899_) );
	INVX1 INVX1_879 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_6900_) );
	OAI22X1 OAI22X1_187 ( .A(_6899_), .B(_6514_), .C(_6563_), .D(_6900_), .Y(_6901_) );
	INVX1 INVX1_880 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_6902_) );
	NAND2X1 NAND2X1_1408 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_6615_), .Y(_6903_) );
	OAI21X1 OAI21X1_231 ( .A(_6902_), .B(_6520_), .C(_6903_), .Y(_6904_) );
	NOR2X1 NOR2X1_814 ( .A(_6901_), .B(_6904_), .Y(_6905_) );
	NAND3X1 NAND3X1_341 ( .A(_6897_), .B(_6898_), .C(_6905_), .Y(_6906_) );
	AND2X2 AND2X2_152 ( .A(_6528_), .B(_6462_), .Y(_6907_) );
	AOI22X1 AOI22X1_1099 ( .A(_6467_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_6907_), .Y(_6908_) );
	AND2X2 AND2X2_153 ( .A(_6526_), .B(_6491_), .Y(_6909_) );
	AND2X2 AND2X2_154 ( .A(_6534_), .B(_6491_), .Y(_6910_) );
	AOI22X1 AOI22X1_1100 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_6910_), .C(_6909_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_6911_) );
	NAND2X1 NAND2X1_1409 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_6619_), .Y(_6912_) );
	NAND2X1 NAND2X1_1410 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_6592_), .Y(_6913_) );
	NAND2X1 NAND2X1_1411 ( .A(_6912_), .B(_6913_), .Y(_6914_) );
	INVX1 INVX1_881 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_6915_) );
	NAND2X1 NAND2X1_1412 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_6591_), .Y(_6916_) );
	OAI21X1 OAI21X1_232 ( .A(_6915_), .B(_6544_), .C(_6916_), .Y(_6917_) );
	NOR2X1 NOR2X1_815 ( .A(_6914_), .B(_6917_), .Y(_6918_) );
	NAND3X1 NAND3X1_342 ( .A(_6908_), .B(_6911_), .C(_6918_), .Y(_6919_) );
	NOR3X1 NOR3X1_584 ( .A(_6906_), .B(_6896_), .C(_6919_), .Y(_6920_) );
	INVX1 INVX1_882 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_6921_) );
	NAND2X1 NAND2X1_1413 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_6507_), .Y(_6922_) );
	OAI21X1 OAI21X1_233 ( .A(_6512_), .B(_6921_), .C(_6922_), .Y(_6923_) );
	AOI21X1 AOI21X1_166 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_6487_), .C(_6923_), .Y(_6924_) );
	INVX1 INVX1_883 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_6925_) );
	INVX1 INVX1_884 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_6926_) );
	OAI22X1 OAI22X1_188 ( .A(_6831_), .B(_6926_), .C(_6925_), .D(_6482_), .Y(_6927_) );
	INVX1 INVX1_885 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_6928_) );
	NAND2X1 NAND2X1_1414 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_6627_), .Y(_6929_) );
	OAI21X1 OAI21X1_234 ( .A(_6492_), .B(_6928_), .C(_6929_), .Y(_6930_) );
	NOR2X1 NOR2X1_816 ( .A(_6930_), .B(_6927_), .Y(_6931_) );
	INVX1 INVX1_886 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_6932_) );
	INVX1 INVX1_887 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_6933_) );
	OAI22X1 OAI22X1_189 ( .A(_6579_), .B(_6933_), .C(_6932_), .D(_6580_), .Y(_6934_) );
	INVX1 INVX1_888 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_6935_) );
	NAND2X1 NAND2X1_1415 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_6626_), .Y(_6936_) );
	OAI21X1 OAI21X1_235 ( .A(_6935_), .B(_6562_), .C(_6936_), .Y(_6937_) );
	NOR2X1 NOR2X1_817 ( .A(_6937_), .B(_6934_), .Y(_6938_) );
	NAND3X1 NAND3X1_343 ( .A(_6924_), .B(_6938_), .C(_6931_), .Y(_6939_) );
	AOI22X1 AOI22X1_1101 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_6584_), .C(_6585_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_6940_) );
	AOI22X1 AOI22X1_1102 ( .A(_6587_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_6588_), .Y(_6941_) );
	NAND2X1 NAND2X1_1416 ( .A(_6940_), .B(_6941_), .Y(_6942_) );
	AOI22X1 AOI22X1_1103 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_6595_), .C(_6594_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_6943_) );
	AOI22X1 AOI22X1_1104 ( .A(_6538_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_6545_), .Y(_6944_) );
	NAND2X1 NAND2X1_1417 ( .A(_6943_), .B(_6944_), .Y(_6945_) );
	NOR2X1 NOR2X1_818 ( .A(_6942_), .B(_6945_), .Y(_6946_) );
	AOI22X1 AOI22X1_1105 ( .A(_6599_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_6600_), .Y(_6947_) );
	AOI22X1 AOI22X1_1106 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_6835_), .C(_6602_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_6948_) );
	NAND2X1 NAND2X1_1418 ( .A(_6948_), .B(_6947_), .Y(_6949_) );
	AOI22X1 AOI22X1_1107 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_6606_), .C(_6607_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_6950_) );
	AOI22X1 AOI22X1_1108 ( .A(_6609_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_6610_), .Y(_6951_) );
	NAND2X1 NAND2X1_1419 ( .A(_6951_), .B(_6950_), .Y(_6952_) );
	NOR2X1 NOR2X1_819 ( .A(_6949_), .B(_6952_), .Y(_6953_) );
	NAND2X1 NAND2X1_1420 ( .A(_6953_), .B(_6946_), .Y(_6954_) );
	AOI22X1 AOI22X1_1109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_6616_), .C(_6517_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_6955_) );
	AOI22X1 AOI22X1_1110 ( .A(_6540_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_6618_), .Y(_6956_) );
	NAND2X1 NAND2X1_1421 ( .A(_6955_), .B(_6956_), .Y(_6957_) );
	AOI22X1 AOI22X1_1111 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_6624_), .C(_6622_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_6958_) );
	AOI22X1 AOI22X1_1112 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_6554_), .C(_6603_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_6959_) );
	NAND2X1 NAND2X1_1422 ( .A(_6959_), .B(_6958_), .Y(_6960_) );
	NOR2X1 NOR2X1_820 ( .A(_6960_), .B(_6957_), .Y(_6961_) );
	AOI22X1 AOI22X1_1113 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_6631_), .C(_6632_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_6962_) );
	NAND2X1 NAND2X1_1423 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_6634_), .Y(_6963_) );
	NAND2X1 NAND2X1_1424 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_6636_), .Y(_6964_) );
	NAND3X1 NAND3X1_344 ( .A(_6963_), .B(_6964_), .C(_6962_), .Y(_6965_) );
	AOI22X1 AOI22X1_1114 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_6640_), .C(_6639_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_6966_) );
	AOI22X1 AOI22X1_1115 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_6643_), .C(_6642_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_6967_) );
	NAND2X1 NAND2X1_1425 ( .A(_6966_), .B(_6967_), .Y(_6968_) );
	NOR2X1 NOR2X1_821 ( .A(_6968_), .B(_6965_), .Y(_6969_) );
	NAND2X1 NAND2X1_1426 ( .A(_6961_), .B(_6969_), .Y(_6970_) );
	NOR3X1 NOR3X1_585 ( .A(_6954_), .B(_6939_), .C(_6970_), .Y(_6971_) );
	NAND2X1 NAND2X1_1427 ( .A(wData[59]), .B(_6673_), .Y(_6972_) );
	OAI21X1 OAI21X1_236 ( .A(_6457_), .B(wBusy_bF_buf2), .C(_6972_), .Y(_6973_) );
	NAND2X1 NAND2X1_1428 ( .A(wData[7]), .B(_6664_), .Y(_6974_) );
	NAND2X1 NAND2X1_1429 ( .A(wData[55]), .B(_6674_), .Y(_6975_) );
	AOI22X1 AOI22X1_1116 ( .A(wData[63]), .B(_6676_), .C(_6666_), .D(wData[31]), .Y(_6976_) );
	NAND3X1 NAND3X1_345 ( .A(_6974_), .B(_6975_), .C(_6976_), .Y(_6977_) );
	OR2X2 OR2X2_78 ( .A(_6977_), .B(_6973_), .Y(_6978_) );
	INVX1 INVX1_889 ( .A(wData[51]), .Y(_6979_) );
	NAND2X1 NAND2X1_1430 ( .A(wData[47]), .B(_6677_), .Y(_6980_) );
	OAI21X1 OAI21X1_237 ( .A(_6979_), .B(_6689_), .C(_6980_), .Y(_6981_) );
	AOI21X1 AOI21X1_167 ( .A(wData[3]), .B(_6684_), .C(_6981_), .Y(_6982_) );
	AOI22X1 AOI22X1_1117 ( .A(_6690_), .B(wData[11]), .C(wData[15]), .D(_6691_), .Y(_6983_) );
	AOI22X1 AOI22X1_1118 ( .A(_6653_), .B(wData[23]), .C(wData[27]), .D(_6660_), .Y(_6984_) );
	AND2X2 AND2X2_155 ( .A(_6983_), .B(_6984_), .Y(_6985_) );
	NAND2X1 NAND2X1_1431 ( .A(wData[39]), .B(_6682_), .Y(_6986_) );
	NAND2X1 NAND2X1_1432 ( .A(wData[43]), .B(_6680_), .Y(_6987_) );
	NAND2X1 NAND2X1_1433 ( .A(_6986_), .B(_6987_), .Y(_6988_) );
	NAND2X1 NAND2X1_1434 ( .A(wData[19]), .B(_6656_), .Y(_6989_) );
	NAND2X1 NAND2X1_1435 ( .A(wData[35]), .B(_6670_), .Y(_6990_) );
	NAND2X1 NAND2X1_1436 ( .A(_6989_), .B(_6990_), .Y(_6991_) );
	NOR2X1 NOR2X1_822 ( .A(_6988_), .B(_6991_), .Y(_6992_) );
	NAND3X1 NAND3X1_346 ( .A(_6985_), .B(_6982_), .C(_6992_), .Y(_6993_) );
	NOR2X1 NOR2X1_823 ( .A(_6978_), .B(_6993_), .Y(_6994_) );
	AOI21X1 AOI21X1_168 ( .A(_6920_), .B(_6971_), .C(_6994_), .Y(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_3_) );
	INVX1 INVX1_890 ( .A(wSelec[143]), .Y(_6995_) );
	NOR2X1 NOR2X1_824 ( .A(wBusy_bF_buf1), .B(_6995_), .Y(_6996_) );
	INVX1 INVX1_891 ( .A(_6996_), .Y(_6997_) );
	INVX1 INVX1_892 ( .A(wSelec[153]), .Y(_6998_) );
	NAND2X1 NAND2X1_1437 ( .A(wSelec[152]), .B(_6998_), .Y(_6999_) );
	INVX2 INVX2_23 ( .A(_6999_), .Y(_7000_) );
	OR2X2 OR2X2_79 ( .A(wSelec[149]), .B(wSelec[148]), .Y(_7001_) );
	INVX1 INVX1_893 ( .A(wSelec[151]), .Y(_7002_) );
	NAND2X1 NAND2X1_1438 ( .A(wSelec[150]), .B(_7002_), .Y(_7003_) );
	NOR2X1 NOR2X1_825 ( .A(_7001_), .B(_7003_), .Y(_7004_) );
	AND2X2 AND2X2_156 ( .A(_7004_), .B(_7000_), .Y(_7005_) );
	AOI21X1 AOI21X1_169 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_7005_), .C(_6997_), .Y(_7006_) );
	INVX1 INVX1_894 ( .A(wSelec[149]), .Y(_7007_) );
	NAND2X1 NAND2X1_1439 ( .A(wSelec[148]), .B(_7007_), .Y(_7008_) );
	OR2X2 OR2X2_80 ( .A(wSelec[150]), .B(wSelec[151]), .Y(_7009_) );
	NOR2X1 NOR2X1_826 ( .A(_7009_), .B(_7008_), .Y(_7010_) );
	NAND2X1 NAND2X1_1440 ( .A(_7000_), .B(_7010_), .Y(_7011_) );
	INVX1 INVX1_895 ( .A(_7011_), .Y(_7012_) );
	INVX1 INVX1_896 ( .A(wSelec[148]), .Y(_7013_) );
	NAND2X1 NAND2X1_1441 ( .A(wSelec[149]), .B(_7013_), .Y(_7014_) );
	INVX1 INVX1_897 ( .A(wSelec[150]), .Y(_7015_) );
	NAND2X1 NAND2X1_1442 ( .A(wSelec[151]), .B(_7015_), .Y(_7016_) );
	NOR2X1 NOR2X1_827 ( .A(_7014_), .B(_7016_), .Y(_7017_) );
	NAND2X1 NAND2X1_1443 ( .A(wSelec[152]), .B(wSelec[153]), .Y(_7018_) );
	INVX1 INVX1_898 ( .A(_7018_), .Y(_7019_) );
	NAND2X1 NAND2X1_1444 ( .A(_7019_), .B(_7017_), .Y(_7020_) );
	INVX1 INVX1_899 ( .A(_7020_), .Y(_7021_) );
	AOI22X1 AOI22X1_1119 ( .A(_7012_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_7021_), .Y(_7022_) );
	OR2X2 OR2X2_81 ( .A(_7008_), .B(_7009_), .Y(_7023_) );
	OR2X2 OR2X2_82 ( .A(wSelec[152]), .B(wSelec[153]), .Y(_7024_) );
	NOR2X1 NOR2X1_828 ( .A(_7024_), .B(_7023_), .Y(_7025_) );
	NOR2X1 NOR2X1_829 ( .A(_7003_), .B(_7008_), .Y(_7026_) );
	INVX1 INVX1_900 ( .A(wSelec[152]), .Y(_7027_) );
	NAND2X1 NAND2X1_1445 ( .A(wSelec[153]), .B(_7027_), .Y(_7028_) );
	INVX2 INVX2_24 ( .A(_7028_), .Y(_7029_) );
	NAND2X1 NAND2X1_1446 ( .A(_7029_), .B(_7026_), .Y(_7030_) );
	INVX1 INVX1_901 ( .A(_7030_), .Y(_7031_) );
	AOI22X1 AOI22X1_1120 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_7025_), .C(_7031_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_7032_) );
	NAND3X1 NAND3X1_347 ( .A(_7006_), .B(_7032_), .C(_7022_), .Y(_7033_) );
	NOR2X1 NOR2X1_830 ( .A(wSelec[149]), .B(wSelec[148]), .Y(_7034_) );
	NOR2X1 NOR2X1_831 ( .A(wSelec[150]), .B(wSelec[151]), .Y(_7035_) );
	NAND2X1 NAND2X1_1447 ( .A(_7034_), .B(_7035_), .Y(_7036_) );
	NOR2X1 NOR2X1_832 ( .A(_6999_), .B(_7036_), .Y(_7037_) );
	NAND2X1 NAND2X1_1448 ( .A(wSelec[149]), .B(wSelec[148]), .Y(_7038_) );
	NOR3X1 NOR3X1_586 ( .A(_7009_), .B(_7038_), .C(_6999_), .Y(_7039_) );
	AOI22X1 AOI22X1_1121 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_7039_), .C(_7037_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_7040_) );
	INVX1 INVX1_902 ( .A(_7024_), .Y(_7041_) );
	NOR2X1 NOR2X1_833 ( .A(_7009_), .B(_7014_), .Y(_7042_) );
	AND2X2 AND2X2_157 ( .A(_7042_), .B(_7041_), .Y(_7043_) );
	NAND2X1 NAND2X1_1449 ( .A(wSelec[150]), .B(wSelec[151]), .Y(_7044_) );
	NOR3X1 NOR3X1_587 ( .A(_7018_), .B(_7038_), .C(_7044_), .Y(_7045_) );
	AOI22X1 AOI22X1_1122 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_7045_), .C(_7043_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_7046_) );
	INVX1 INVX1_903 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_7047_) );
	INVX1 INVX1_904 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_7048_) );
	NOR2X1 NOR2X1_834 ( .A(_7008_), .B(_7016_), .Y(_7049_) );
	NAND2X1 NAND2X1_1450 ( .A(_7019_), .B(_7049_), .Y(_7050_) );
	NOR2X1 NOR2X1_835 ( .A(_7038_), .B(_7044_), .Y(_7051_) );
	NAND2X1 NAND2X1_1451 ( .A(_7051_), .B(_7029_), .Y(_7052_) );
	OAI22X1 OAI22X1_190 ( .A(_7047_), .B(_7052_), .C(_7050_), .D(_7048_), .Y(_7053_) );
	INVX1 INVX1_905 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_7054_) );
	NOR3X1 NOR3X1_588 ( .A(_6999_), .B(_7014_), .C(_7016_), .Y(_7055_) );
	NAND2X1 NAND2X1_1452 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_7055_), .Y(_7056_) );
	NOR2X1 NOR2X1_836 ( .A(_7038_), .B(_7003_), .Y(_7057_) );
	NAND2X1 NAND2X1_1453 ( .A(_7029_), .B(_7057_), .Y(_7058_) );
	OAI21X1 OAI21X1_238 ( .A(_7054_), .B(_7058_), .C(_7056_), .Y(_7059_) );
	NOR2X1 NOR2X1_837 ( .A(_7053_), .B(_7059_), .Y(_7060_) );
	NAND3X1 NAND3X1_348 ( .A(_7040_), .B(_7046_), .C(_7060_), .Y(_7061_) );
	INVX1 INVX1_906 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_7062_) );
	INVX1 INVX1_907 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_7063_) );
	NOR2X1 NOR2X1_838 ( .A(_7003_), .B(_7014_), .Y(_7064_) );
	NAND2X1 NAND2X1_1454 ( .A(_7000_), .B(_7064_), .Y(_7065_) );
	NOR2X1 NOR2X1_839 ( .A(_7001_), .B(_7016_), .Y(_7066_) );
	NAND2X1 NAND2X1_1455 ( .A(_7000_), .B(_7066_), .Y(_7067_) );
	OAI22X1 OAI22X1_191 ( .A(_7067_), .B(_7062_), .C(_7063_), .D(_7065_), .Y(_7068_) );
	INVX1 INVX1_908 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_7069_) );
	INVX1 INVX1_909 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_7070_) );
	NAND2X1 NAND2X1_1456 ( .A(_7029_), .B(_7064_), .Y(_7071_) );
	NOR2X1 NOR2X1_840 ( .A(_7038_), .B(_7009_), .Y(_7072_) );
	NAND2X1 NAND2X1_1457 ( .A(_7029_), .B(_7072_), .Y(_7073_) );
	OAI22X1 OAI22X1_192 ( .A(_7069_), .B(_7073_), .C(_7071_), .D(_7070_), .Y(_7074_) );
	NOR2X1 NOR2X1_841 ( .A(_7074_), .B(_7068_), .Y(_7075_) );
	NOR3X1 NOR3X1_589 ( .A(_7008_), .B(_7044_), .C(_7028_), .Y(_7076_) );
	NAND2X1 NAND2X1_1458 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_7076_), .Y(_7077_) );
	NOR3X1 NOR3X1_590 ( .A(_7016_), .B(_7038_), .C(_7028_), .Y(_7078_) );
	NAND2X1 NAND2X1_1459 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_7078_), .Y(_7079_) );
	NAND2X1 NAND2X1_1460 ( .A(_7077_), .B(_7079_), .Y(_7080_) );
	INVX1 INVX1_910 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_7081_) );
	NAND2X1 NAND2X1_1461 ( .A(_7019_), .B(_7004_), .Y(_7082_) );
	NOR3X1 NOR3X1_591 ( .A(_7014_), .B(_7016_), .C(_7028_), .Y(_7083_) );
	NAND2X1 NAND2X1_1462 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_7083_), .Y(_7084_) );
	OAI21X1 OAI21X1_239 ( .A(_7081_), .B(_7082_), .C(_7084_), .Y(_7085_) );
	NOR2X1 NOR2X1_842 ( .A(_7080_), .B(_7085_), .Y(_7086_) );
	NAND2X1 NAND2X1_1463 ( .A(_7075_), .B(_7086_), .Y(_7087_) );
	NOR3X1 NOR3X1_592 ( .A(_7033_), .B(_7087_), .C(_7061_), .Y(_7088_) );
	NAND2X1 NAND2X1_1464 ( .A(_7000_), .B(_7057_), .Y(_7089_) );
	INVX1 INVX1_911 ( .A(_7089_), .Y(_7090_) );
	INVX1 INVX1_912 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_7091_) );
	NOR3X1 NOR3X1_593 ( .A(_7001_), .B(_7024_), .C(_7003_), .Y(_7092_) );
	NAND2X1 NAND2X1_1465 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_7092_), .Y(_7093_) );
	NAND2X1 NAND2X1_1466 ( .A(_7041_), .B(_7064_), .Y(_7094_) );
	OAI21X1 OAI21X1_240 ( .A(_7094_), .B(_7091_), .C(_7093_), .Y(_7095_) );
	AOI21X1 AOI21X1_170 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_7090_), .C(_7095_), .Y(_7096_) );
	INVX1 INVX1_913 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_7097_) );
	INVX1 INVX1_914 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_7098_) );
	NOR2X1 NOR2X1_843 ( .A(_7044_), .B(_7001_), .Y(_7099_) );
	NAND2X1 NAND2X1_1467 ( .A(_7000_), .B(_7099_), .Y(_7100_) );
	NAND2X1 NAND2X1_1468 ( .A(_7041_), .B(_7026_), .Y(_7101_) );
	OAI22X1 OAI22X1_193 ( .A(_7098_), .B(_7100_), .C(_7101_), .D(_7097_), .Y(_7102_) );
	INVX1 INVX1_915 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_7103_) );
	INVX1 INVX1_916 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_7104_) );
	NAND2X1 NAND2X1_1469 ( .A(_7000_), .B(_7026_), .Y(_7105_) );
	NAND2X1 NAND2X1_1470 ( .A(_7041_), .B(_7072_), .Y(_7106_) );
	OAI22X1 OAI22X1_194 ( .A(_7103_), .B(_7106_), .C(_7105_), .D(_7104_), .Y(_7107_) );
	NOR2X1 NOR2X1_844 ( .A(_7102_), .B(_7107_), .Y(_7108_) );
	INVX1 INVX1_917 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_7109_) );
	NOR3X1 NOR3X1_594 ( .A(_7024_), .B(_7038_), .C(_7003_), .Y(_7110_) );
	NAND2X1 NAND2X1_1471 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_7110_), .Y(_7111_) );
	OR2X2 OR2X2_83 ( .A(_7036_), .B(_7018_), .Y(_7112_) );
	OAI21X1 OAI21X1_241 ( .A(_7109_), .B(_7112_), .C(_7111_), .Y(_7113_) );
	INVX1 INVX1_918 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_7114_) );
	INVX1 INVX1_919 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_7115_) );
	NOR2X1 NOR2X1_845 ( .A(_7044_), .B(_7014_), .Y(_7116_) );
	NAND2X1 NAND2X1_1472 ( .A(_7000_), .B(_7116_), .Y(_7117_) );
	NAND2X1 NAND2X1_1473 ( .A(_7019_), .B(_7010_), .Y(_7118_) );
	OAI22X1 OAI22X1_195 ( .A(_7117_), .B(_7115_), .C(_7114_), .D(_7118_), .Y(_7119_) );
	NOR2X1 NOR2X1_846 ( .A(_7113_), .B(_7119_), .Y(_7120_) );
	NAND3X1 NAND3X1_349 ( .A(_7096_), .B(_7120_), .C(_7108_), .Y(_7121_) );
	NOR3X1 NOR3X1_595 ( .A(_7001_), .B(_7009_), .C(_7024_), .Y(_7122_) );
	NOR3X1 NOR3X1_596 ( .A(_7018_), .B(_7044_), .C(_7008_), .Y(_7123_) );
	AOI22X1 AOI22X1_1123 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_7122_), .C(_7123_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_7124_) );
	NOR3X1 NOR3X1_597 ( .A(_7018_), .B(_7044_), .C(_7014_), .Y(_7125_) );
	NOR3X1 NOR3X1_598 ( .A(_7018_), .B(_7038_), .C(_7016_), .Y(_7126_) );
	AOI22X1 AOI22X1_1124 ( .A(_7125_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_7126_), .Y(_7127_) );
	NAND2X1 NAND2X1_1474 ( .A(_7124_), .B(_7127_), .Y(_7128_) );
	NOR3X1 NOR3X1_599 ( .A(_7016_), .B(_7001_), .C(_7028_), .Y(_7129_) );
	NOR3X1 NOR3X1_600 ( .A(_7008_), .B(_7016_), .C(_7028_), .Y(_7130_) );
	AOI22X1 AOI22X1_1125 ( .A(_7129_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_7130_), .Y(_7131_) );
	NOR3X1 NOR3X1_601 ( .A(_6999_), .B(_7044_), .C(_7008_), .Y(_7132_) );
	NOR3X1 NOR3X1_602 ( .A(_7038_), .B(_7044_), .C(_6999_), .Y(_7133_) );
	AOI22X1 AOI22X1_1126 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_7133_), .C(_7132_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_7134_) );
	NAND2X1 NAND2X1_1475 ( .A(_7134_), .B(_7131_), .Y(_7135_) );
	NOR2X1 NOR2X1_847 ( .A(_7128_), .B(_7135_), .Y(_7136_) );
	NOR3X1 NOR3X1_603 ( .A(_7024_), .B(_7044_), .C(_7008_), .Y(_7137_) );
	NOR3X1 NOR3X1_604 ( .A(_7024_), .B(_7044_), .C(_7014_), .Y(_7138_) );
	AOI22X1 AOI22X1_1127 ( .A(_7137_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_7138_), .Y(_7139_) );
	NOR3X1 NOR3X1_605 ( .A(_7024_), .B(_7038_), .C(_7016_), .Y(_7140_) );
	NOR3X1 NOR3X1_606 ( .A(_6999_), .B(_7009_), .C(_7014_), .Y(_7141_) );
	AOI22X1 AOI22X1_1128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_7140_), .C(_7141_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_7142_) );
	NAND2X1 NAND2X1_1476 ( .A(_7139_), .B(_7142_), .Y(_7143_) );
	NOR3X1 NOR3X1_607 ( .A(_7038_), .B(_7044_), .C(_7024_), .Y(_7144_) );
	NOR3X1 NOR3X1_608 ( .A(_7014_), .B(_7009_), .C(_7028_), .Y(_7145_) );
	AOI22X1 AOI22X1_1129 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_7144_), .C(_7145_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_7146_) );
	NOR3X1 NOR3X1_609 ( .A(_7001_), .B(_7009_), .C(_7028_), .Y(_7147_) );
	NOR3X1 NOR3X1_610 ( .A(_7001_), .B(_7044_), .C(_7028_), .Y(_7148_) );
	AOI22X1 AOI22X1_1130 ( .A(_7147_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_7148_), .Y(_7149_) );
	NAND2X1 NAND2X1_1477 ( .A(_7149_), .B(_7146_), .Y(_7150_) );
	NOR2X1 NOR2X1_848 ( .A(_7143_), .B(_7150_), .Y(_7151_) );
	NAND2X1 NAND2X1_1478 ( .A(_7151_), .B(_7136_), .Y(_7152_) );
	NOR3X1 NOR3X1_611 ( .A(_6999_), .B(_7038_), .C(_7016_), .Y(_7153_) );
	NOR3X1 NOR3X1_612 ( .A(_7009_), .B(_7018_), .C(_7014_), .Y(_7154_) );
	AOI22X1 AOI22X1_1131 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_7154_), .C(_7153_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_7155_) );
	NOR3X1 NOR3X1_613 ( .A(_7003_), .B(_7001_), .C(_7028_), .Y(_7156_) );
	NOR3X1 NOR3X1_614 ( .A(_7014_), .B(_7044_), .C(_7028_), .Y(_7157_) );
	AOI22X1 AOI22X1_1132 ( .A(_7156_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_7157_), .Y(_7158_) );
	NAND2X1 NAND2X1_1479 ( .A(_7155_), .B(_7158_), .Y(_7159_) );
	NOR3X1 NOR3X1_615 ( .A(_6999_), .B(_7008_), .C(_7016_), .Y(_7160_) );
	NAND2X1 NAND2X1_1480 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_7160_), .Y(_7161_) );
	NOR3X1 NOR3X1_616 ( .A(_7018_), .B(_7038_), .C(_7003_), .Y(_7162_) );
	NAND2X1 NAND2X1_1481 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_7162_), .Y(_7163_) );
	NOR3X1 NOR3X1_617 ( .A(_7001_), .B(_7044_), .C(_7024_), .Y(_7164_) );
	NOR3X1 NOR3X1_618 ( .A(_7001_), .B(_7018_), .C(_7016_), .Y(_7165_) );
	AOI22X1 AOI22X1_1133 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_7164_), .C(_7165_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_7166_) );
	NAND3X1 NAND3X1_350 ( .A(_7161_), .B(_7163_), .C(_7166_), .Y(_7167_) );
	NOR2X1 NOR2X1_849 ( .A(_7167_), .B(_7159_), .Y(_7168_) );
	NOR3X1 NOR3X1_619 ( .A(_7001_), .B(_7024_), .C(_7016_), .Y(_7169_) );
	NOR3X1 NOR3X1_620 ( .A(_7003_), .B(_7018_), .C(_7008_), .Y(_7170_) );
	AOI22X1 AOI22X1_1134 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_7169_), .C(_7170_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_7171_) );
	NOR3X1 NOR3X1_621 ( .A(_7003_), .B(_7018_), .C(_7014_), .Y(_7172_) );
	NAND2X1 NAND2X1_1482 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_7172_), .Y(_7173_) );
	NOR3X1 NOR3X1_622 ( .A(_7008_), .B(_7009_), .C(_7028_), .Y(_7174_) );
	NAND2X1 NAND2X1_1483 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_7174_), .Y(_7175_) );
	NAND3X1 NAND3X1_351 ( .A(_7173_), .B(_7175_), .C(_7171_), .Y(_7176_) );
	NOR3X1 NOR3X1_623 ( .A(_7008_), .B(_7024_), .C(_7016_), .Y(_7177_) );
	NOR3X1 NOR3X1_624 ( .A(_7018_), .B(_7044_), .C(_7001_), .Y(_7178_) );
	AOI22X1 AOI22X1_1135 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_7178_), .C(_7177_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_7179_) );
	NOR3X1 NOR3X1_625 ( .A(_7014_), .B(_7024_), .C(_7016_), .Y(_7180_) );
	NOR3X1 NOR3X1_626 ( .A(_7018_), .B(_7038_), .C(_7009_), .Y(_7181_) );
	AOI22X1 AOI22X1_1136 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_7181_), .C(_7180_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_7182_) );
	NAND2X1 NAND2X1_1484 ( .A(_7179_), .B(_7182_), .Y(_7183_) );
	NOR2X1 NOR2X1_850 ( .A(_7183_), .B(_7176_), .Y(_7184_) );
	NAND2X1 NAND2X1_1485 ( .A(_7168_), .B(_7184_), .Y(_7185_) );
	NOR3X1 NOR3X1_627 ( .A(_7152_), .B(_7121_), .C(_7185_), .Y(_7186_) );
	INVX1 INVX1_920 ( .A(wSelec[145]), .Y(_7187_) );
	NAND2X1 NAND2X1_1486 ( .A(wSelec[144]), .B(_7187_), .Y(_7188_) );
	INVX1 INVX1_921 ( .A(wSelec[147]), .Y(_7189_) );
	NAND2X1 NAND2X1_1487 ( .A(wSelec[146]), .B(_7189_), .Y(_7190_) );
	NOR2X1 NOR2X1_851 ( .A(_7188_), .B(_7190_), .Y(_7191_) );
	NOR2X1 NOR2X1_852 ( .A(wSelec[145]), .B(wSelec[144]), .Y(_7192_) );
	INVX1 INVX1_922 ( .A(_7192_), .Y(_7193_) );
	NOR2X1 NOR2X1_853 ( .A(_7190_), .B(_7193_), .Y(_7194_) );
	AOI22X1 AOI22X1_1137 ( .A(wData[20]), .B(_7191_), .C(_7194_), .D(wData[16]), .Y(_7195_) );
	INVX1 INVX1_923 ( .A(wSelec[144]), .Y(_7196_) );
	NAND2X1 NAND2X1_1488 ( .A(wSelec[145]), .B(_7196_), .Y(_7197_) );
	NOR2X1 NOR2X1_854 ( .A(_7197_), .B(_7190_), .Y(_7198_) );
	NAND2X1 NAND2X1_1489 ( .A(wData[24]), .B(_7198_), .Y(_7199_) );
	INVX1 INVX1_924 ( .A(wSelec[146]), .Y(_7200_) );
	NAND2X1 NAND2X1_1490 ( .A(_7200_), .B(_7189_), .Y(_7201_) );
	NOR2X1 NOR2X1_855 ( .A(_7188_), .B(_7201_), .Y(_7202_) );
	NAND2X1 NAND2X1_1491 ( .A(wSelec[145]), .B(wSelec[144]), .Y(_7203_) );
	NOR2X1 NOR2X1_856 ( .A(_7203_), .B(_7190_), .Y(_7204_) );
	AOI22X1 AOI22X1_1138 ( .A(_7204_), .B(wData[28]), .C(wData[4]), .D(_7202_), .Y(_7205_) );
	NAND3X1 NAND3X1_352 ( .A(_7199_), .B(_7205_), .C(_7195_), .Y(_7206_) );
	NAND2X1 NAND2X1_1492 ( .A(wSelec[147]), .B(_7200_), .Y(_7207_) );
	NOR2X1 NOR2X1_857 ( .A(_7207_), .B(_7193_), .Y(_7208_) );
	NAND2X1 NAND2X1_1493 ( .A(wData[32]), .B(_7208_), .Y(_7209_) );
	NAND2X1 NAND2X1_1494 ( .A(wSelec[146]), .B(wSelec[147]), .Y(_7210_) );
	NOR2X1 NOR2X1_858 ( .A(_7210_), .B(_7197_), .Y(_7211_) );
	NOR2X1 NOR2X1_859 ( .A(_7210_), .B(_7188_), .Y(_7212_) );
	AOI22X1 AOI22X1_1139 ( .A(_7211_), .B(wData[56]), .C(wData[52]), .D(_7212_), .Y(_7213_) );
	NOR2X1 NOR2X1_860 ( .A(_7203_), .B(_7210_), .Y(_7214_) );
	NOR2X1 NOR2X1_861 ( .A(_7203_), .B(_7207_), .Y(_7215_) );
	AOI22X1 AOI22X1_1140 ( .A(wData[60]), .B(_7214_), .C(_7215_), .D(wData[44]), .Y(_7216_) );
	NAND3X1 NAND3X1_353 ( .A(_7209_), .B(_7216_), .C(_7213_), .Y(_7217_) );
	NOR2X1 NOR2X1_862 ( .A(_7197_), .B(_7207_), .Y(_7218_) );
	NAND2X1 NAND2X1_1495 ( .A(wData[40]), .B(_7218_), .Y(_7219_) );
	NOR2X1 NOR2X1_863 ( .A(_7207_), .B(_7188_), .Y(_7220_) );
	NAND2X1 NAND2X1_1496 ( .A(wData[36]), .B(_7220_), .Y(_7221_) );
	NOR2X1 NOR2X1_864 ( .A(_7201_), .B(_7193_), .Y(_7222_) );
	NAND2X1 NAND2X1_1497 ( .A(wData[0]), .B(_7222_), .Y(_7223_) );
	NAND3X1 NAND3X1_354 ( .A(_7219_), .B(_7221_), .C(_7223_), .Y(_7224_) );
	INVX1 INVX1_925 ( .A(wData[48]), .Y(_7225_) );
	NOR2X1 NOR2X1_865 ( .A(_7200_), .B(_7189_), .Y(_7226_) );
	NAND2X1 NAND2X1_1498 ( .A(_7192_), .B(_7226_), .Y(_7227_) );
	NOR2X1 NOR2X1_866 ( .A(_7197_), .B(_7201_), .Y(_7228_) );
	NOR2X1 NOR2X1_867 ( .A(_7203_), .B(_7201_), .Y(_7229_) );
	AOI22X1 AOI22X1_1141 ( .A(_7228_), .B(wData[8]), .C(wData[12]), .D(_7229_), .Y(_7230_) );
	OAI21X1 OAI21X1_242 ( .A(_7225_), .B(_7227_), .C(_7230_), .Y(_7231_) );
	OR2X2 OR2X2_84 ( .A(_7231_), .B(_7224_), .Y(_7232_) );
	NOR3X1 NOR3X1_628 ( .A(_7206_), .B(_7217_), .C(_7232_), .Y(_7233_) );
	AND2X2 AND2X2_158 ( .A(_7233_), .B(_6997_), .Y(_7234_) );
	AOI21X1 AOI21X1_171 ( .A(_7088_), .B(_7186_), .C(_7234_), .Y(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_0_) );
	INVX1 INVX1_926 ( .A(_7105_), .Y(_7235_) );
	AOI21X1 AOI21X1_172 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_7235_), .C(_6997_), .Y(_7236_) );
	AOI22X1 AOI22X1_1142 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_7005_), .C(_7021_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_7237_) );
	AOI22X1 AOI22X1_1143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_7025_), .C(_7031_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_7238_) );
	NAND3X1 NAND3X1_355 ( .A(_7236_), .B(_7237_), .C(_7238_), .Y(_7239_) );
	INVX1 INVX1_927 ( .A(_7065_), .Y(_7240_) );
	AOI22X1 AOI22X1_1144 ( .A(_7090_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_7240_), .Y(_7241_) );
	AOI22X1 AOI22X1_1145 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_7164_), .C(_7043_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_7242_) );
	INVX1 INVX1_928 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_7243_) );
	INVX1 INVX1_929 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_7244_) );
	OAI22X1 OAI22X1_196 ( .A(_7243_), .B(_7052_), .C(_7050_), .D(_7244_), .Y(_7245_) );
	INVX1 INVX1_930 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_7246_) );
	NAND2X1 NAND2X1_1499 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_7153_), .Y(_7247_) );
	OAI21X1 OAI21X1_243 ( .A(_7246_), .B(_7058_), .C(_7247_), .Y(_7248_) );
	NOR2X1 NOR2X1_868 ( .A(_7245_), .B(_7248_), .Y(_7249_) );
	NAND3X1 NAND3X1_356 ( .A(_7241_), .B(_7242_), .C(_7249_), .Y(_7250_) );
	INVX1 INVX1_931 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_7251_) );
	NAND2X1 NAND2X1_1500 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_7037_), .Y(_7252_) );
	OAI21X1 OAI21X1_244 ( .A(_7251_), .B(_7067_), .C(_7252_), .Y(_7253_) );
	INVX1 INVX1_932 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_7254_) );
	INVX1 INVX1_933 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_7255_) );
	OAI22X1 OAI22X1_197 ( .A(_7254_), .B(_7073_), .C(_7071_), .D(_7255_), .Y(_7256_) );
	NOR2X1 NOR2X1_869 ( .A(_7256_), .B(_7253_), .Y(_7257_) );
	AOI22X1 AOI22X1_1146 ( .A(_7157_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_7130_), .Y(_7258_) );
	AND2X2 AND2X2_159 ( .A(_7004_), .B(_7019_), .Y(_7259_) );
	AOI22X1 AOI22X1_1147 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_7129_), .C(_7259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_7260_) );
	NAND3X1 NAND3X1_357 ( .A(_7258_), .B(_7260_), .C(_7257_), .Y(_7261_) );
	NOR3X1 NOR3X1_629 ( .A(_7261_), .B(_7239_), .C(_7250_), .Y(_7262_) );
	INVX1 INVX1_934 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_7263_) );
	NAND2X1 NAND2X1_1501 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_7092_), .Y(_7264_) );
	OAI21X1 OAI21X1_245 ( .A(_7094_), .B(_7263_), .C(_7264_), .Y(_7265_) );
	AOI21X1 AOI21X1_173 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_7141_), .C(_7265_), .Y(_7266_) );
	INVX1 INVX1_935 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_7267_) );
	INVX1 INVX1_936 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_7268_) );
	OAI22X1 OAI22X1_198 ( .A(_7268_), .B(_7100_), .C(_7101_), .D(_7267_), .Y(_7269_) );
	INVX1 INVX1_937 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_7270_) );
	NAND2X1 NAND2X1_1502 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_7110_), .Y(_7271_) );
	OAI21X1 OAI21X1_246 ( .A(_7011_), .B(_7270_), .C(_7271_), .Y(_7272_) );
	NOR2X1 NOR2X1_870 ( .A(_7272_), .B(_7269_), .Y(_7273_) );
	INVX1 INVX1_938 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_7274_) );
	INVX1 INVX1_939 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_7275_) );
	OAI22X1 OAI22X1_199 ( .A(_7106_), .B(_7275_), .C(_7112_), .D(_7274_), .Y(_7276_) );
	INVX1 INVX1_940 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_7277_) );
	NOR2X1 NOR2X1_871 ( .A(_7277_), .B(_7117_), .Y(_7278_) );
	INVX1 INVX1_941 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_7279_) );
	NOR2X1 NOR2X1_872 ( .A(_7279_), .B(_7118_), .Y(_7280_) );
	NOR3X1 NOR3X1_630 ( .A(_7278_), .B(_7276_), .C(_7280_), .Y(_7281_) );
	NAND3X1 NAND3X1_358 ( .A(_7273_), .B(_7266_), .C(_7281_), .Y(_7282_) );
	AOI22X1 AOI22X1_1148 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_7122_), .C(_7123_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_7283_) );
	AOI22X1 AOI22X1_1149 ( .A(_7125_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_7126_), .Y(_7284_) );
	NAND2X1 NAND2X1_1503 ( .A(_7283_), .B(_7284_), .Y(_7285_) );
	AOI22X1 AOI22X1_1150 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_7133_), .C(_7132_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_7286_) );
	AOI22X1 AOI22X1_1151 ( .A(_7076_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_7083_), .Y(_7287_) );
	NAND2X1 NAND2X1_1504 ( .A(_7286_), .B(_7287_), .Y(_7288_) );
	NOR2X1 NOR2X1_873 ( .A(_7285_), .B(_7288_), .Y(_7289_) );
	AOI22X1 AOI22X1_1152 ( .A(_7137_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_7138_), .Y(_7290_) );
	AOI22X1 AOI22X1_1153 ( .A(_7039_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_7140_), .Y(_7291_) );
	NAND2X1 NAND2X1_1505 ( .A(_7290_), .B(_7291_), .Y(_7292_) );
	AOI22X1 AOI22X1_1154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_7144_), .C(_7145_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_7293_) );
	AOI22X1 AOI22X1_1155 ( .A(_7147_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_7148_), .Y(_7294_) );
	NAND2X1 NAND2X1_1506 ( .A(_7294_), .B(_7293_), .Y(_7295_) );
	NOR2X1 NOR2X1_874 ( .A(_7292_), .B(_7295_), .Y(_7296_) );
	NAND2X1 NAND2X1_1507 ( .A(_7296_), .B(_7289_), .Y(_7297_) );
	AOI22X1 AOI22X1_1156 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_7154_), .C(_7055_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_7298_) );
	AOI22X1 AOI22X1_1157 ( .A(_7078_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_7156_), .Y(_7299_) );
	NAND2X1 NAND2X1_1508 ( .A(_7298_), .B(_7299_), .Y(_7300_) );
	AOI22X1 AOI22X1_1158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_7045_), .C(_7165_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_7301_) );
	NAND2X1 NAND2X1_1509 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_7160_), .Y(_7302_) );
	NAND2X1 NAND2X1_1510 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_7162_), .Y(_7303_) );
	NAND3X1 NAND3X1_359 ( .A(_7302_), .B(_7303_), .C(_7301_), .Y(_7304_) );
	NOR2X1 NOR2X1_875 ( .A(_7304_), .B(_7300_), .Y(_7305_) );
	AOI22X1 AOI22X1_1159 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_7169_), .C(_7170_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_7306_) );
	NAND2X1 NAND2X1_1511 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_7172_), .Y(_7307_) );
	NAND2X1 NAND2X1_1512 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_7174_), .Y(_7308_) );
	NAND3X1 NAND3X1_360 ( .A(_7307_), .B(_7308_), .C(_7306_), .Y(_7309_) );
	AOI22X1 AOI22X1_1160 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_7178_), .C(_7177_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_7310_) );
	AOI22X1 AOI22X1_1161 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_7181_), .C(_7180_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_7311_) );
	NAND2X1 NAND2X1_1513 ( .A(_7310_), .B(_7311_), .Y(_7312_) );
	NOR2X1 NOR2X1_876 ( .A(_7312_), .B(_7309_), .Y(_7313_) );
	NAND2X1 NAND2X1_1514 ( .A(_7305_), .B(_7313_), .Y(_7314_) );
	NOR3X1 NOR3X1_631 ( .A(_7297_), .B(_7282_), .C(_7314_), .Y(_7315_) );
	AOI21X1 AOI21X1_174 ( .A(wData[21]), .B(_7191_), .C(_6996_), .Y(_7316_) );
	AOI22X1 AOI22X1_1162 ( .A(_7194_), .B(wData[17]), .C(wData[1]), .D(_7222_), .Y(_7317_) );
	AOI22X1 AOI22X1_1163 ( .A(_7215_), .B(wData[45]), .C(wData[25]), .D(_7198_), .Y(_7318_) );
	NAND3X1 NAND3X1_361 ( .A(_7316_), .B(_7318_), .C(_7317_), .Y(_7319_) );
	NAND3X1 NAND3X1_362 ( .A(wData[49]), .B(_7192_), .C(_7226_), .Y(_7320_) );
	AOI22X1 AOI22X1_1164 ( .A(wData[61]), .B(_7214_), .C(_7202_), .D(wData[5]), .Y(_7321_) );
	AND2X2 AND2X2_160 ( .A(_7321_), .B(_7320_), .Y(_7322_) );
	AOI22X1 AOI22X1_1165 ( .A(_7211_), .B(wData[57]), .C(wData[41]), .D(_7218_), .Y(_7323_) );
	AOI22X1 AOI22X1_1166 ( .A(wData[53]), .B(_7212_), .C(_7208_), .D(wData[33]), .Y(_7324_) );
	AND2X2 AND2X2_161 ( .A(_7324_), .B(_7323_), .Y(_7325_) );
	AOI22X1 AOI22X1_1167 ( .A(_7228_), .B(wData[9]), .C(wData[13]), .D(_7229_), .Y(_7326_) );
	AOI22X1 AOI22X1_1168 ( .A(_7204_), .B(wData[29]), .C(wData[37]), .D(_7220_), .Y(_7327_) );
	AND2X2 AND2X2_162 ( .A(_7326_), .B(_7327_), .Y(_7328_) );
	NAND3X1 NAND3X1_363 ( .A(_7322_), .B(_7328_), .C(_7325_), .Y(_7329_) );
	NOR2X1 NOR2X1_877 ( .A(_7319_), .B(_7329_), .Y(_7330_) );
	AOI21X1 AOI21X1_175 ( .A(_7262_), .B(_7315_), .C(_7330_), .Y(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_1_) );
	AOI21X1 AOI21X1_176 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_7235_), .C(_6997_), .Y(_7331_) );
	INVX1 INVX1_942 ( .A(_7094_), .Y(_7332_) );
	AOI22X1 AOI22X1_1169 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_7005_), .C(_7332_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_7333_) );
	INVX1 INVX1_943 ( .A(_7106_), .Y(_7334_) );
	AOI22X1 AOI22X1_1170 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_7141_), .C(_7334_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_7335_) );
	NAND3X1 NAND3X1_364 ( .A(_7335_), .B(_7331_), .C(_7333_), .Y(_7336_) );
	AOI22X1 AOI22X1_1171 ( .A(_7090_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_7240_), .Y(_7337_) );
	AOI22X1 AOI22X1_1172 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_7039_), .C(_7012_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_7338_) );
	INVX1 INVX1_944 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_7339_) );
	NAND2X1 NAND2X1_1515 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_7129_), .Y(_7340_) );
	OAI21X1 OAI21X1_247 ( .A(_7339_), .B(_7101_), .C(_7340_), .Y(_7341_) );
	INVX1 INVX1_945 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_7342_) );
	NAND2X1 NAND2X1_1516 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_7055_), .Y(_7343_) );
	OAI21X1 OAI21X1_248 ( .A(_7342_), .B(_7058_), .C(_7343_), .Y(_7344_) );
	NOR2X1 NOR2X1_878 ( .A(_7341_), .B(_7344_), .Y(_7345_) );
	NAND3X1 NAND3X1_365 ( .A(_7337_), .B(_7338_), .C(_7345_), .Y(_7346_) );
	INVX1 INVX1_946 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_7347_) );
	NAND2X1 NAND2X1_1517 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_7037_), .Y(_7348_) );
	OAI21X1 OAI21X1_249 ( .A(_7347_), .B(_7067_), .C(_7348_), .Y(_7349_) );
	INVX1 INVX1_947 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_7350_) );
	INVX1 INVX1_948 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_7351_) );
	OAI22X1 OAI22X1_200 ( .A(_7350_), .B(_7073_), .C(_7071_), .D(_7351_), .Y(_7352_) );
	NOR2X1 NOR2X1_879 ( .A(_7352_), .B(_7349_), .Y(_7353_) );
	AOI22X1 AOI22X1_1173 ( .A(_7157_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_7130_), .Y(_7354_) );
	AND2X2 AND2X2_163 ( .A(_7029_), .B(_7051_), .Y(_7355_) );
	AOI22X1 AOI22X1_1174 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_7355_), .C(_7259_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_7356_) );
	NAND3X1 NAND3X1_366 ( .A(_7354_), .B(_7356_), .C(_7353_), .Y(_7357_) );
	NOR3X1 NOR3X1_632 ( .A(_7357_), .B(_7336_), .C(_7346_), .Y(_7358_) );
	INVX1 INVX1_949 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_7359_) );
	NOR3X1 NOR3X1_633 ( .A(_7359_), .B(_7024_), .C(_7023_), .Y(_7360_) );
	AND2X2 AND2X2_164 ( .A(_7045_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_7361_) );
	AND2X2 AND2X2_165 ( .A(_7165_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_7362_) );
	NOR3X1 NOR3X1_634 ( .A(_7362_), .B(_7361_), .C(_7360_), .Y(_7363_) );
	INVX1 INVX1_950 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_7364_) );
	INVX1 INVX1_951 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_7365_) );
	OAI22X1 OAI22X1_201 ( .A(_7365_), .B(_7100_), .C(_7050_), .D(_7364_), .Y(_7366_) );
	INVX1 INVX1_952 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_7367_) );
	INVX1 INVX1_953 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_7368_) );
	NAND2X1 NAND2X1_1518 ( .A(_7041_), .B(_7042_), .Y(_7369_) );
	OAI22X1 OAI22X1_202 ( .A(_7369_), .B(_7368_), .C(_7367_), .D(_7020_), .Y(_7370_) );
	NOR2X1 NOR2X1_880 ( .A(_7366_), .B(_7370_), .Y(_7371_) );
	INVX1 INVX1_954 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_7372_) );
	NOR3X1 NOR3X1_635 ( .A(_7001_), .B(_7018_), .C(_7009_), .Y(_7373_) );
	NAND2X1 NAND2X1_1519 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_7373_), .Y(_7374_) );
	OAI21X1 OAI21X1_250 ( .A(_7030_), .B(_7372_), .C(_7374_), .Y(_7375_) );
	INVX1 INVX1_955 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_7376_) );
	INVX1 INVX1_956 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_7377_) );
	OAI22X1 OAI22X1_203 ( .A(_7117_), .B(_7377_), .C(_7376_), .D(_7118_), .Y(_7378_) );
	NOR2X1 NOR2X1_881 ( .A(_7375_), .B(_7378_), .Y(_7379_) );
	NAND3X1 NAND3X1_367 ( .A(_7363_), .B(_7379_), .C(_7371_), .Y(_7380_) );
	AOI22X1 AOI22X1_1175 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_7122_), .C(_7123_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_7381_) );
	AOI22X1 AOI22X1_1176 ( .A(_7125_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_7126_), .Y(_7382_) );
	NAND2X1 NAND2X1_1520 ( .A(_7381_), .B(_7382_), .Y(_7383_) );
	AOI22X1 AOI22X1_1177 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_7133_), .C(_7132_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_7384_) );
	AOI22X1 AOI22X1_1178 ( .A(_7076_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_7083_), .Y(_7385_) );
	NAND2X1 NAND2X1_1521 ( .A(_7384_), .B(_7385_), .Y(_7386_) );
	NOR2X1 NOR2X1_882 ( .A(_7383_), .B(_7386_), .Y(_7387_) );
	AOI22X1 AOI22X1_1179 ( .A(_7137_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_7138_), .Y(_7388_) );
	AOI22X1 AOI22X1_1180 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_7164_), .C(_7140_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_7389_) );
	NAND2X1 NAND2X1_1522 ( .A(_7389_), .B(_7388_), .Y(_7390_) );
	AOI22X1 AOI22X1_1181 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_7144_), .C(_7145_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_7391_) );
	AOI22X1 AOI22X1_1182 ( .A(_7147_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_7148_), .Y(_7392_) );
	NAND2X1 NAND2X1_1523 ( .A(_7392_), .B(_7391_), .Y(_7393_) );
	NOR2X1 NOR2X1_883 ( .A(_7390_), .B(_7393_), .Y(_7394_) );
	NAND2X1 NAND2X1_1524 ( .A(_7394_), .B(_7387_), .Y(_7395_) );
	AOI22X1 AOI22X1_1183 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_7154_), .C(_7153_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_7396_) );
	AOI22X1 AOI22X1_1184 ( .A(_7078_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_7156_), .Y(_7397_) );
	NAND2X1 NAND2X1_1525 ( .A(_7396_), .B(_7397_), .Y(_7398_) );
	AOI22X1 AOI22X1_1185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_7162_), .C(_7160_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_7399_) );
	AOI22X1 AOI22X1_1186 ( .A(_7092_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_7110_), .Y(_7400_) );
	NAND2X1 NAND2X1_1526 ( .A(_7400_), .B(_7399_), .Y(_7401_) );
	NOR2X1 NOR2X1_884 ( .A(_7401_), .B(_7398_), .Y(_7402_) );
	AOI22X1 AOI22X1_1187 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_7169_), .C(_7170_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_7403_) );
	NAND2X1 NAND2X1_1527 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_7172_), .Y(_7404_) );
	NAND2X1 NAND2X1_1528 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_7174_), .Y(_7405_) );
	NAND3X1 NAND3X1_368 ( .A(_7404_), .B(_7405_), .C(_7403_), .Y(_7406_) );
	AOI22X1 AOI22X1_1188 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_7178_), .C(_7177_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_7407_) );
	AOI22X1 AOI22X1_1189 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_7181_), .C(_7180_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_7408_) );
	NAND2X1 NAND2X1_1529 ( .A(_7407_), .B(_7408_), .Y(_7409_) );
	NOR2X1 NOR2X1_885 ( .A(_7409_), .B(_7406_), .Y(_7410_) );
	NAND2X1 NAND2X1_1530 ( .A(_7402_), .B(_7410_), .Y(_7411_) );
	NOR3X1 NOR3X1_636 ( .A(_7395_), .B(_7380_), .C(_7411_), .Y(_7412_) );
	AOI22X1 AOI22X1_1190 ( .A(_7218_), .B(wData[42]), .C(wData[38]), .D(_7220_), .Y(_7413_) );
	AOI22X1 AOI22X1_1191 ( .A(_7215_), .B(wData[46]), .C(_7222_), .D(wData[2]), .Y(_7414_) );
	NAND2X1 NAND2X1_1531 ( .A(_7413_), .B(_7414_), .Y(_7415_) );
	AOI21X1 AOI21X1_177 ( .A(wData[34]), .B(_7208_), .C(_7415_), .Y(_7416_) );
	INVX1 INVX1_957 ( .A(wData[50]), .Y(_7417_) );
	AOI22X1 AOI22X1_1192 ( .A(_7228_), .B(wData[10]), .C(wData[14]), .D(_7229_), .Y(_7418_) );
	OAI21X1 OAI21X1_251 ( .A(_7417_), .B(_7227_), .C(_7418_), .Y(_7419_) );
	AOI22X1 AOI22X1_1193 ( .A(_7191_), .B(wData[22]), .C(wData[18]), .D(_7194_), .Y(_7420_) );
	NAND2X1 NAND2X1_1532 ( .A(wData[26]), .B(_7198_), .Y(_7421_) );
	AOI22X1 AOI22X1_1194 ( .A(_7204_), .B(wData[30]), .C(wData[6]), .D(_7202_), .Y(_7422_) );
	NAND3X1 NAND3X1_369 ( .A(_7421_), .B(_7422_), .C(_7420_), .Y(_7423_) );
	NOR2X1 NOR2X1_886 ( .A(_7419_), .B(_7423_), .Y(_7424_) );
	NAND2X1 NAND2X1_1533 ( .A(wData[58]), .B(_7211_), .Y(_7425_) );
	NAND2X1 NAND2X1_1534 ( .A(wData[54]), .B(_7212_), .Y(_7426_) );
	NAND2X1 NAND2X1_1535 ( .A(_7425_), .B(_7426_), .Y(_7427_) );
	AOI21X1 AOI21X1_178 ( .A(wData[62]), .B(_7214_), .C(_7427_), .Y(_7428_) );
	NAND3X1 NAND3X1_370 ( .A(_7416_), .B(_7428_), .C(_7424_), .Y(_7429_) );
	NOR2X1 NOR2X1_887 ( .A(_6996_), .B(_7429_), .Y(_7430_) );
	AOI21X1 AOI21X1_179 ( .A(_7358_), .B(_7412_), .C(_7430_), .Y(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_2_) );
	AOI21X1 AOI21X1_180 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_7240_), .C(_6997_), .Y(_7431_) );
	AOI22X1 AOI22X1_1195 ( .A(_7012_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_7332_), .Y(_7432_) );
	AOI22X1 AOI22X1_1196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_7334_), .C(_7090_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_7433_) );
	NAND3X1 NAND3X1_371 ( .A(_7433_), .B(_7431_), .C(_7432_), .Y(_7434_) );
	AOI22X1 AOI22X1_1197 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_7039_), .C(_7037_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_7435_) );
	AOI22X1 AOI22X1_1198 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_7110_), .C(_7235_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_7436_) );
	INVX1 INVX1_958 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_7437_) );
	INVX1 INVX1_959 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_7438_) );
	OAI22X1 OAI22X1_204 ( .A(_7437_), .B(_7052_), .C(_7101_), .D(_7438_), .Y(_7439_) );
	INVX1 INVX1_960 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_7440_) );
	NAND2X1 NAND2X1_1536 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_7153_), .Y(_7441_) );
	OAI21X1 OAI21X1_252 ( .A(_7440_), .B(_7058_), .C(_7441_), .Y(_7442_) );
	NOR2X1 NOR2X1_888 ( .A(_7439_), .B(_7442_), .Y(_7443_) );
	NAND3X1 NAND3X1_372 ( .A(_7435_), .B(_7436_), .C(_7443_), .Y(_7444_) );
	AND2X2 AND2X2_166 ( .A(_7066_), .B(_7000_), .Y(_7445_) );
	AOI22X1 AOI22X1_1199 ( .A(_7005_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_7445_), .Y(_7446_) );
	AND2X2 AND2X2_167 ( .A(_7064_), .B(_7029_), .Y(_7447_) );
	AND2X2 AND2X2_168 ( .A(_7072_), .B(_7029_), .Y(_7448_) );
	AOI22X1 AOI22X1_1200 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_7448_), .C(_7447_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_7449_) );
	NAND2X1 NAND2X1_1537 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_7157_), .Y(_7450_) );
	NAND2X1 NAND2X1_1538 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_7130_), .Y(_7451_) );
	NAND2X1 NAND2X1_1539 ( .A(_7450_), .B(_7451_), .Y(_7452_) );
	INVX1 INVX1_961 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_7453_) );
	NAND2X1 NAND2X1_1540 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_7129_), .Y(_7454_) );
	OAI21X1 OAI21X1_253 ( .A(_7453_), .B(_7082_), .C(_7454_), .Y(_7455_) );
	NOR2X1 NOR2X1_889 ( .A(_7452_), .B(_7455_), .Y(_7456_) );
	NAND3X1 NAND3X1_373 ( .A(_7446_), .B(_7449_), .C(_7456_), .Y(_7457_) );
	NOR3X1 NOR3X1_637 ( .A(_7444_), .B(_7434_), .C(_7457_), .Y(_7458_) );
	INVX1 INVX1_962 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_7459_) );
	NAND2X1 NAND2X1_1541 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_7045_), .Y(_7460_) );
	OAI21X1 OAI21X1_254 ( .A(_7050_), .B(_7459_), .C(_7460_), .Y(_7461_) );
	AOI21X1 AOI21X1_181 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_7025_), .C(_7461_), .Y(_7462_) );
	INVX1 INVX1_963 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_7463_) );
	INVX1 INVX1_964 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_7464_) );
	OAI22X1 OAI22X1_205 ( .A(_7369_), .B(_7464_), .C(_7463_), .D(_7020_), .Y(_7465_) );
	INVX1 INVX1_965 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_7466_) );
	NAND2X1 NAND2X1_1542 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_7165_), .Y(_7467_) );
	OAI21X1 OAI21X1_255 ( .A(_7030_), .B(_7466_), .C(_7467_), .Y(_7468_) );
	NOR2X1 NOR2X1_890 ( .A(_7468_), .B(_7465_), .Y(_7469_) );
	INVX1 INVX1_966 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_7470_) );
	INVX1 INVX1_967 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_7471_) );
	OAI22X1 OAI22X1_206 ( .A(_7117_), .B(_7471_), .C(_7470_), .D(_7118_), .Y(_7472_) );
	INVX1 INVX1_968 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_7473_) );
	NAND2X1 NAND2X1_1543 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_7164_), .Y(_7474_) );
	OAI21X1 OAI21X1_256 ( .A(_7473_), .B(_7100_), .C(_7474_), .Y(_7475_) );
	NOR2X1 NOR2X1_891 ( .A(_7475_), .B(_7472_), .Y(_7476_) );
	NAND3X1 NAND3X1_374 ( .A(_7462_), .B(_7476_), .C(_7469_), .Y(_7477_) );
	AOI22X1 AOI22X1_1201 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_7122_), .C(_7123_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_7478_) );
	AOI22X1 AOI22X1_1202 ( .A(_7125_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_7126_), .Y(_7479_) );
	NAND2X1 NAND2X1_1544 ( .A(_7478_), .B(_7479_), .Y(_7480_) );
	AOI22X1 AOI22X1_1203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_7133_), .C(_7132_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_7481_) );
	AOI22X1 AOI22X1_1204 ( .A(_7076_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_7083_), .Y(_7482_) );
	NAND2X1 NAND2X1_1545 ( .A(_7481_), .B(_7482_), .Y(_7483_) );
	NOR2X1 NOR2X1_892 ( .A(_7480_), .B(_7483_), .Y(_7484_) );
	AOI22X1 AOI22X1_1205 ( .A(_7137_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_7138_), .Y(_7485_) );
	AOI22X1 AOI22X1_1206 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_7373_), .C(_7140_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_7486_) );
	NAND2X1 NAND2X1_1546 ( .A(_7486_), .B(_7485_), .Y(_7487_) );
	AOI22X1 AOI22X1_1207 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_7144_), .C(_7145_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_7488_) );
	AOI22X1 AOI22X1_1208 ( .A(_7147_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_7148_), .Y(_7489_) );
	NAND2X1 NAND2X1_1547 ( .A(_7489_), .B(_7488_), .Y(_7490_) );
	NOR2X1 NOR2X1_893 ( .A(_7487_), .B(_7490_), .Y(_7491_) );
	NAND2X1 NAND2X1_1548 ( .A(_7491_), .B(_7484_), .Y(_7492_) );
	AOI22X1 AOI22X1_1209 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_7154_), .C(_7055_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_7493_) );
	AOI22X1 AOI22X1_1210 ( .A(_7078_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_7156_), .Y(_7494_) );
	NAND2X1 NAND2X1_1549 ( .A(_7493_), .B(_7494_), .Y(_7495_) );
	AOI22X1 AOI22X1_1211 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_7162_), .C(_7160_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_7496_) );
	AOI22X1 AOI22X1_1212 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_7092_), .C(_7141_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_7497_) );
	NAND2X1 NAND2X1_1550 ( .A(_7497_), .B(_7496_), .Y(_7498_) );
	NOR2X1 NOR2X1_894 ( .A(_7498_), .B(_7495_), .Y(_7499_) );
	AOI22X1 AOI22X1_1213 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_7169_), .C(_7170_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_7500_) );
	NAND2X1 NAND2X1_1551 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_7172_), .Y(_7501_) );
	NAND2X1 NAND2X1_1552 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_7174_), .Y(_7502_) );
	NAND3X1 NAND3X1_375 ( .A(_7501_), .B(_7502_), .C(_7500_), .Y(_7503_) );
	AOI22X1 AOI22X1_1214 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_7178_), .C(_7177_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_7504_) );
	AOI22X1 AOI22X1_1215 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_7181_), .C(_7180_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_7505_) );
	NAND2X1 NAND2X1_1553 ( .A(_7504_), .B(_7505_), .Y(_7506_) );
	NOR2X1 NOR2X1_895 ( .A(_7506_), .B(_7503_), .Y(_7507_) );
	NAND2X1 NAND2X1_1554 ( .A(_7499_), .B(_7507_), .Y(_7508_) );
	NOR3X1 NOR3X1_638 ( .A(_7492_), .B(_7477_), .C(_7508_), .Y(_7509_) );
	NAND2X1 NAND2X1_1555 ( .A(wData[59]), .B(_7211_), .Y(_7510_) );
	OAI21X1 OAI21X1_257 ( .A(_6995_), .B(wBusy_bF_buf0), .C(_7510_), .Y(_7511_) );
	NAND2X1 NAND2X1_1556 ( .A(wData[7]), .B(_7202_), .Y(_7512_) );
	NAND2X1 NAND2X1_1557 ( .A(wData[55]), .B(_7212_), .Y(_7513_) );
	AOI22X1 AOI22X1_1216 ( .A(wData[63]), .B(_7214_), .C(_7204_), .D(wData[31]), .Y(_7514_) );
	NAND3X1 NAND3X1_376 ( .A(_7512_), .B(_7513_), .C(_7514_), .Y(_7515_) );
	OR2X2 OR2X2_85 ( .A(_7515_), .B(_7511_), .Y(_7516_) );
	INVX1 INVX1_969 ( .A(wData[51]), .Y(_7517_) );
	NAND2X1 NAND2X1_1558 ( .A(wData[47]), .B(_7215_), .Y(_7518_) );
	OAI21X1 OAI21X1_258 ( .A(_7517_), .B(_7227_), .C(_7518_), .Y(_7519_) );
	AOI21X1 AOI21X1_182 ( .A(wData[3]), .B(_7222_), .C(_7519_), .Y(_7520_) );
	AOI22X1 AOI22X1_1217 ( .A(_7228_), .B(wData[11]), .C(wData[15]), .D(_7229_), .Y(_7521_) );
	AOI22X1 AOI22X1_1218 ( .A(_7191_), .B(wData[23]), .C(wData[27]), .D(_7198_), .Y(_7522_) );
	AND2X2 AND2X2_169 ( .A(_7521_), .B(_7522_), .Y(_7523_) );
	NAND2X1 NAND2X1_1559 ( .A(wData[39]), .B(_7220_), .Y(_7524_) );
	NAND2X1 NAND2X1_1560 ( .A(wData[43]), .B(_7218_), .Y(_7525_) );
	NAND2X1 NAND2X1_1561 ( .A(_7524_), .B(_7525_), .Y(_7526_) );
	NAND2X1 NAND2X1_1562 ( .A(wData[19]), .B(_7194_), .Y(_7527_) );
	NAND2X1 NAND2X1_1563 ( .A(wData[35]), .B(_7208_), .Y(_7528_) );
	NAND2X1 NAND2X1_1564 ( .A(_7527_), .B(_7528_), .Y(_7529_) );
	NOR2X1 NOR2X1_896 ( .A(_7526_), .B(_7529_), .Y(_7530_) );
	NAND3X1 NAND3X1_377 ( .A(_7523_), .B(_7520_), .C(_7530_), .Y(_7531_) );
	NOR2X1 NOR2X1_897 ( .A(_7516_), .B(_7531_), .Y(_7532_) );
	AOI21X1 AOI21X1_183 ( .A(_7458_), .B(_7509_), .C(_7532_), .Y(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_3_) );
	INVX1 INVX1_970 ( .A(wSelec[154]), .Y(_7533_) );
	NOR2X1 NOR2X1_898 ( .A(wBusy_bF_buf4), .B(_7533_), .Y(_7534_) );
	INVX1 INVX1_971 ( .A(_7534_), .Y(_7535_) );
	INVX1 INVX1_972 ( .A(wSelec[164]), .Y(_7536_) );
	NAND2X1 NAND2X1_1565 ( .A(wSelec[163]), .B(_7536_), .Y(_7537_) );
	INVX2 INVX2_25 ( .A(_7537_), .Y(_7538_) );
	OR2X2 OR2X2_86 ( .A(wSelec[160]), .B(wSelec[159]), .Y(_7539_) );
	INVX1 INVX1_973 ( .A(wSelec[162]), .Y(_7540_) );
	NAND2X1 NAND2X1_1566 ( .A(wSelec[161]), .B(_7540_), .Y(_7541_) );
	NOR2X1 NOR2X1_899 ( .A(_7539_), .B(_7541_), .Y(_7542_) );
	AND2X2 AND2X2_170 ( .A(_7542_), .B(_7538_), .Y(_7543_) );
	AOI21X1 AOI21X1_184 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_7543_), .C(_7535_), .Y(_7544_) );
	INVX1 INVX1_974 ( .A(wSelec[160]), .Y(_7545_) );
	NAND2X1 NAND2X1_1567 ( .A(wSelec[159]), .B(_7545_), .Y(_7546_) );
	OR2X2 OR2X2_87 ( .A(wSelec[161]), .B(wSelec[162]), .Y(_7547_) );
	NOR2X1 NOR2X1_900 ( .A(_7547_), .B(_7546_), .Y(_7548_) );
	NAND2X1 NAND2X1_1568 ( .A(_7538_), .B(_7548_), .Y(_7549_) );
	INVX1 INVX1_975 ( .A(_7549_), .Y(_7550_) );
	INVX1 INVX1_976 ( .A(wSelec[159]), .Y(_7551_) );
	NAND2X1 NAND2X1_1569 ( .A(wSelec[160]), .B(_7551_), .Y(_7552_) );
	INVX1 INVX1_977 ( .A(wSelec[161]), .Y(_7553_) );
	NAND2X1 NAND2X1_1570 ( .A(wSelec[162]), .B(_7553_), .Y(_7554_) );
	NOR2X1 NOR2X1_901 ( .A(_7552_), .B(_7554_), .Y(_7555_) );
	NAND2X1 NAND2X1_1571 ( .A(wSelec[163]), .B(wSelec[164]), .Y(_7556_) );
	INVX1 INVX1_978 ( .A(_7556_), .Y(_7557_) );
	NAND2X1 NAND2X1_1572 ( .A(_7557_), .B(_7555_), .Y(_7558_) );
	INVX1 INVX1_979 ( .A(_7558_), .Y(_7559_) );
	AOI22X1 AOI22X1_1219 ( .A(_7550_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_7559_), .Y(_7560_) );
	OR2X2 OR2X2_88 ( .A(_7546_), .B(_7547_), .Y(_7561_) );
	OR2X2 OR2X2_89 ( .A(wSelec[163]), .B(wSelec[164]), .Y(_7562_) );
	NOR2X1 NOR2X1_902 ( .A(_7562_), .B(_7561_), .Y(_7563_) );
	NOR2X1 NOR2X1_903 ( .A(_7541_), .B(_7546_), .Y(_7564_) );
	INVX1 INVX1_980 ( .A(wSelec[163]), .Y(_7565_) );
	NAND2X1 NAND2X1_1573 ( .A(wSelec[164]), .B(_7565_), .Y(_7566_) );
	INVX2 INVX2_26 ( .A(_7566_), .Y(_7567_) );
	NAND2X1 NAND2X1_1574 ( .A(_7567_), .B(_7564_), .Y(_7568_) );
	INVX1 INVX1_981 ( .A(_7568_), .Y(_7569_) );
	AOI22X1 AOI22X1_1220 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_7563_), .C(_7569_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_7570_) );
	NAND3X1 NAND3X1_378 ( .A(_7544_), .B(_7570_), .C(_7560_), .Y(_7571_) );
	NOR2X1 NOR2X1_904 ( .A(wSelec[160]), .B(wSelec[159]), .Y(_7572_) );
	NOR2X1 NOR2X1_905 ( .A(wSelec[161]), .B(wSelec[162]), .Y(_7573_) );
	NAND2X1 NAND2X1_1575 ( .A(_7572_), .B(_7573_), .Y(_7574_) );
	NOR2X1 NOR2X1_906 ( .A(_7537_), .B(_7574_), .Y(_7575_) );
	NAND2X1 NAND2X1_1576 ( .A(wSelec[160]), .B(wSelec[159]), .Y(_7576_) );
	NOR3X1 NOR3X1_639 ( .A(_7547_), .B(_7576_), .C(_7537_), .Y(_7577_) );
	AOI22X1 AOI22X1_1221 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_7577_), .C(_7575_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_7578_) );
	INVX1 INVX1_982 ( .A(_7562_), .Y(_7579_) );
	NOR2X1 NOR2X1_907 ( .A(_7547_), .B(_7552_), .Y(_7580_) );
	AND2X2 AND2X2_171 ( .A(_7580_), .B(_7579_), .Y(_7581_) );
	NAND2X1 NAND2X1_1577 ( .A(wSelec[161]), .B(wSelec[162]), .Y(_7582_) );
	NOR3X1 NOR3X1_640 ( .A(_7556_), .B(_7576_), .C(_7582_), .Y(_7583_) );
	AOI22X1 AOI22X1_1222 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_7583_), .C(_7581_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_7584_) );
	INVX1 INVX1_983 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_7585_) );
	INVX1 INVX1_984 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_7586_) );
	NOR2X1 NOR2X1_908 ( .A(_7546_), .B(_7554_), .Y(_7587_) );
	NAND2X1 NAND2X1_1578 ( .A(_7557_), .B(_7587_), .Y(_7588_) );
	NOR2X1 NOR2X1_909 ( .A(_7576_), .B(_7582_), .Y(_7589_) );
	NAND2X1 NAND2X1_1579 ( .A(_7589_), .B(_7567_), .Y(_7590_) );
	OAI22X1 OAI22X1_207 ( .A(_7585_), .B(_7590_), .C(_7588_), .D(_7586_), .Y(_7591_) );
	INVX1 INVX1_985 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_7592_) );
	NOR3X1 NOR3X1_641 ( .A(_7537_), .B(_7552_), .C(_7554_), .Y(_7593_) );
	NAND2X1 NAND2X1_1580 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_7593_), .Y(_7594_) );
	NOR2X1 NOR2X1_910 ( .A(_7576_), .B(_7541_), .Y(_7595_) );
	NAND2X1 NAND2X1_1581 ( .A(_7567_), .B(_7595_), .Y(_7596_) );
	OAI21X1 OAI21X1_259 ( .A(_7592_), .B(_7596_), .C(_7594_), .Y(_7597_) );
	NOR2X1 NOR2X1_911 ( .A(_7591_), .B(_7597_), .Y(_7598_) );
	NAND3X1 NAND3X1_379 ( .A(_7578_), .B(_7584_), .C(_7598_), .Y(_7599_) );
	INVX1 INVX1_986 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_7600_) );
	INVX1 INVX1_987 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_7601_) );
	NOR2X1 NOR2X1_912 ( .A(_7541_), .B(_7552_), .Y(_7602_) );
	NAND2X1 NAND2X1_1582 ( .A(_7538_), .B(_7602_), .Y(_7603_) );
	NOR2X1 NOR2X1_913 ( .A(_7539_), .B(_7554_), .Y(_7604_) );
	NAND2X1 NAND2X1_1583 ( .A(_7538_), .B(_7604_), .Y(_7605_) );
	OAI22X1 OAI22X1_208 ( .A(_7605_), .B(_7600_), .C(_7601_), .D(_7603_), .Y(_7606_) );
	INVX1 INVX1_988 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_7607_) );
	INVX1 INVX1_989 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_7608_) );
	NAND2X1 NAND2X1_1584 ( .A(_7567_), .B(_7602_), .Y(_7609_) );
	NOR2X1 NOR2X1_914 ( .A(_7576_), .B(_7547_), .Y(_7610_) );
	NAND2X1 NAND2X1_1585 ( .A(_7567_), .B(_7610_), .Y(_7611_) );
	OAI22X1 OAI22X1_209 ( .A(_7607_), .B(_7611_), .C(_7609_), .D(_7608_), .Y(_7612_) );
	NOR2X1 NOR2X1_915 ( .A(_7612_), .B(_7606_), .Y(_7613_) );
	NOR3X1 NOR3X1_642 ( .A(_7546_), .B(_7582_), .C(_7566_), .Y(_7614_) );
	NAND2X1 NAND2X1_1586 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_7614_), .Y(_7615_) );
	NOR3X1 NOR3X1_643 ( .A(_7554_), .B(_7576_), .C(_7566_), .Y(_7616_) );
	NAND2X1 NAND2X1_1587 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_7616_), .Y(_7617_) );
	NAND2X1 NAND2X1_1588 ( .A(_7615_), .B(_7617_), .Y(_7618_) );
	INVX1 INVX1_990 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_7619_) );
	NAND2X1 NAND2X1_1589 ( .A(_7557_), .B(_7542_), .Y(_7620_) );
	NOR3X1 NOR3X1_644 ( .A(_7552_), .B(_7554_), .C(_7566_), .Y(_7621_) );
	NAND2X1 NAND2X1_1590 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_7621_), .Y(_7622_) );
	OAI21X1 OAI21X1_260 ( .A(_7619_), .B(_7620_), .C(_7622_), .Y(_7623_) );
	NOR2X1 NOR2X1_916 ( .A(_7618_), .B(_7623_), .Y(_7624_) );
	NAND2X1 NAND2X1_1591 ( .A(_7613_), .B(_7624_), .Y(_7625_) );
	NOR3X1 NOR3X1_645 ( .A(_7571_), .B(_7625_), .C(_7599_), .Y(_7626_) );
	NAND2X1 NAND2X1_1592 ( .A(_7538_), .B(_7595_), .Y(_7627_) );
	INVX1 INVX1_991 ( .A(_7627_), .Y(_7628_) );
	INVX1 INVX1_992 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_7629_) );
	NOR3X1 NOR3X1_646 ( .A(_7539_), .B(_7562_), .C(_7541_), .Y(_7630_) );
	NAND2X1 NAND2X1_1593 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_7630_), .Y(_7631_) );
	NAND2X1 NAND2X1_1594 ( .A(_7579_), .B(_7602_), .Y(_7632_) );
	OAI21X1 OAI21X1_261 ( .A(_7632_), .B(_7629_), .C(_7631_), .Y(_7633_) );
	AOI21X1 AOI21X1_185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_7628_), .C(_7633_), .Y(_7634_) );
	INVX1 INVX1_993 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_7635_) );
	INVX1 INVX1_994 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_7636_) );
	NOR2X1 NOR2X1_917 ( .A(_7582_), .B(_7539_), .Y(_7637_) );
	NAND2X1 NAND2X1_1595 ( .A(_7538_), .B(_7637_), .Y(_7638_) );
	NAND2X1 NAND2X1_1596 ( .A(_7579_), .B(_7564_), .Y(_7639_) );
	OAI22X1 OAI22X1_210 ( .A(_7636_), .B(_7638_), .C(_7639_), .D(_7635_), .Y(_7640_) );
	INVX1 INVX1_995 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_7641_) );
	INVX1 INVX1_996 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_7642_) );
	NAND2X1 NAND2X1_1597 ( .A(_7538_), .B(_7564_), .Y(_7643_) );
	NAND2X1 NAND2X1_1598 ( .A(_7579_), .B(_7610_), .Y(_7644_) );
	OAI22X1 OAI22X1_211 ( .A(_7641_), .B(_7644_), .C(_7643_), .D(_7642_), .Y(_7645_) );
	NOR2X1 NOR2X1_918 ( .A(_7640_), .B(_7645_), .Y(_7646_) );
	INVX1 INVX1_997 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_7647_) );
	NOR3X1 NOR3X1_647 ( .A(_7562_), .B(_7576_), .C(_7541_), .Y(_7648_) );
	NAND2X1 NAND2X1_1599 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_7648_), .Y(_7649_) );
	OR2X2 OR2X2_90 ( .A(_7574_), .B(_7556_), .Y(_7650_) );
	OAI21X1 OAI21X1_262 ( .A(_7647_), .B(_7650_), .C(_7649_), .Y(_7651_) );
	INVX1 INVX1_998 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_7652_) );
	INVX1 INVX1_999 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_7653_) );
	NOR2X1 NOR2X1_919 ( .A(_7582_), .B(_7552_), .Y(_7654_) );
	NAND2X1 NAND2X1_1600 ( .A(_7538_), .B(_7654_), .Y(_7655_) );
	NAND2X1 NAND2X1_1601 ( .A(_7557_), .B(_7548_), .Y(_7656_) );
	OAI22X1 OAI22X1_212 ( .A(_7655_), .B(_7653_), .C(_7652_), .D(_7656_), .Y(_7657_) );
	NOR2X1 NOR2X1_920 ( .A(_7651_), .B(_7657_), .Y(_7658_) );
	NAND3X1 NAND3X1_380 ( .A(_7634_), .B(_7658_), .C(_7646_), .Y(_7659_) );
	NOR3X1 NOR3X1_648 ( .A(_7539_), .B(_7547_), .C(_7562_), .Y(_7660_) );
	NOR3X1 NOR3X1_649 ( .A(_7556_), .B(_7582_), .C(_7546_), .Y(_7661_) );
	AOI22X1 AOI22X1_1223 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_7660_), .C(_7661_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_7662_) );
	NOR3X1 NOR3X1_650 ( .A(_7556_), .B(_7582_), .C(_7552_), .Y(_7663_) );
	NOR3X1 NOR3X1_651 ( .A(_7556_), .B(_7576_), .C(_7554_), .Y(_7664_) );
	AOI22X1 AOI22X1_1224 ( .A(_7663_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_7664_), .Y(_7665_) );
	NAND2X1 NAND2X1_1602 ( .A(_7662_), .B(_7665_), .Y(_7666_) );
	NOR3X1 NOR3X1_652 ( .A(_7554_), .B(_7539_), .C(_7566_), .Y(_7667_) );
	NOR3X1 NOR3X1_653 ( .A(_7546_), .B(_7554_), .C(_7566_), .Y(_7668_) );
	AOI22X1 AOI22X1_1225 ( .A(_7667_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_7668_), .Y(_7669_) );
	NOR3X1 NOR3X1_654 ( .A(_7537_), .B(_7582_), .C(_7546_), .Y(_7670_) );
	NOR3X1 NOR3X1_655 ( .A(_7576_), .B(_7582_), .C(_7537_), .Y(_7671_) );
	AOI22X1 AOI22X1_1226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_7671_), .C(_7670_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_7672_) );
	NAND2X1 NAND2X1_1603 ( .A(_7672_), .B(_7669_), .Y(_7673_) );
	NOR2X1 NOR2X1_921 ( .A(_7666_), .B(_7673_), .Y(_7674_) );
	NOR3X1 NOR3X1_656 ( .A(_7562_), .B(_7582_), .C(_7546_), .Y(_7675_) );
	NOR3X1 NOR3X1_657 ( .A(_7562_), .B(_7582_), .C(_7552_), .Y(_7676_) );
	AOI22X1 AOI22X1_1227 ( .A(_7675_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_7676_), .Y(_7677_) );
	NOR3X1 NOR3X1_658 ( .A(_7562_), .B(_7576_), .C(_7554_), .Y(_7678_) );
	NOR3X1 NOR3X1_659 ( .A(_7537_), .B(_7547_), .C(_7552_), .Y(_7679_) );
	AOI22X1 AOI22X1_1228 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_7678_), .C(_7679_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_7680_) );
	NAND2X1 NAND2X1_1604 ( .A(_7677_), .B(_7680_), .Y(_7681_) );
	NOR3X1 NOR3X1_660 ( .A(_7576_), .B(_7582_), .C(_7562_), .Y(_7682_) );
	NOR3X1 NOR3X1_661 ( .A(_7552_), .B(_7547_), .C(_7566_), .Y(_7683_) );
	AOI22X1 AOI22X1_1229 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_7682_), .C(_7683_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_7684_) );
	NOR3X1 NOR3X1_662 ( .A(_7539_), .B(_7547_), .C(_7566_), .Y(_7685_) );
	NOR3X1 NOR3X1_663 ( .A(_7539_), .B(_7582_), .C(_7566_), .Y(_7686_) );
	AOI22X1 AOI22X1_1230 ( .A(_7685_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_7686_), .Y(_7687_) );
	NAND2X1 NAND2X1_1605 ( .A(_7687_), .B(_7684_), .Y(_7688_) );
	NOR2X1 NOR2X1_922 ( .A(_7681_), .B(_7688_), .Y(_7689_) );
	NAND2X1 NAND2X1_1606 ( .A(_7689_), .B(_7674_), .Y(_7690_) );
	NOR3X1 NOR3X1_664 ( .A(_7537_), .B(_7576_), .C(_7554_), .Y(_7691_) );
	NOR3X1 NOR3X1_665 ( .A(_7547_), .B(_7556_), .C(_7552_), .Y(_7692_) );
	AOI22X1 AOI22X1_1231 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_7692_), .C(_7691_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_7693_) );
	NOR3X1 NOR3X1_666 ( .A(_7541_), .B(_7539_), .C(_7566_), .Y(_7694_) );
	NOR3X1 NOR3X1_667 ( .A(_7552_), .B(_7582_), .C(_7566_), .Y(_7695_) );
	AOI22X1 AOI22X1_1232 ( .A(_7694_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_7695_), .Y(_7696_) );
	NAND2X1 NAND2X1_1607 ( .A(_7693_), .B(_7696_), .Y(_7697_) );
	NOR3X1 NOR3X1_668 ( .A(_7537_), .B(_7546_), .C(_7554_), .Y(_7698_) );
	NAND2X1 NAND2X1_1608 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_7698_), .Y(_7699_) );
	NOR3X1 NOR3X1_669 ( .A(_7556_), .B(_7576_), .C(_7541_), .Y(_7700_) );
	NAND2X1 NAND2X1_1609 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_7700_), .Y(_7701_) );
	NOR3X1 NOR3X1_670 ( .A(_7539_), .B(_7582_), .C(_7562_), .Y(_7702_) );
	NOR3X1 NOR3X1_671 ( .A(_7539_), .B(_7556_), .C(_7554_), .Y(_7703_) );
	AOI22X1 AOI22X1_1233 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_7702_), .C(_7703_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_7704_) );
	NAND3X1 NAND3X1_381 ( .A(_7699_), .B(_7701_), .C(_7704_), .Y(_7705_) );
	NOR2X1 NOR2X1_923 ( .A(_7705_), .B(_7697_), .Y(_7706_) );
	NOR3X1 NOR3X1_672 ( .A(_7539_), .B(_7562_), .C(_7554_), .Y(_7707_) );
	NOR3X1 NOR3X1_673 ( .A(_7541_), .B(_7556_), .C(_7546_), .Y(_7708_) );
	AOI22X1 AOI22X1_1234 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_7707_), .C(_7708_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_7709_) );
	NOR3X1 NOR3X1_674 ( .A(_7541_), .B(_7556_), .C(_7552_), .Y(_7710_) );
	NAND2X1 NAND2X1_1610 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_7710_), .Y(_7711_) );
	NOR3X1 NOR3X1_675 ( .A(_7546_), .B(_7547_), .C(_7566_), .Y(_7712_) );
	NAND2X1 NAND2X1_1611 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_7712_), .Y(_7713_) );
	NAND3X1 NAND3X1_382 ( .A(_7711_), .B(_7713_), .C(_7709_), .Y(_7714_) );
	NOR3X1 NOR3X1_676 ( .A(_7546_), .B(_7562_), .C(_7554_), .Y(_7715_) );
	NOR3X1 NOR3X1_677 ( .A(_7556_), .B(_7582_), .C(_7539_), .Y(_7716_) );
	AOI22X1 AOI22X1_1235 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_7716_), .C(_7715_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_7717_) );
	NOR3X1 NOR3X1_678 ( .A(_7552_), .B(_7562_), .C(_7554_), .Y(_7718_) );
	NOR3X1 NOR3X1_679 ( .A(_7556_), .B(_7576_), .C(_7547_), .Y(_7719_) );
	AOI22X1 AOI22X1_1236 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_7719_), .C(_7718_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_7720_) );
	NAND2X1 NAND2X1_1612 ( .A(_7717_), .B(_7720_), .Y(_7721_) );
	NOR2X1 NOR2X1_924 ( .A(_7721_), .B(_7714_), .Y(_7722_) );
	NAND2X1 NAND2X1_1613 ( .A(_7706_), .B(_7722_), .Y(_7723_) );
	NOR3X1 NOR3X1_680 ( .A(_7690_), .B(_7659_), .C(_7723_), .Y(_7724_) );
	INVX1 INVX1_1000 ( .A(wSelec[156]), .Y(_7725_) );
	NAND2X1 NAND2X1_1614 ( .A(wSelec[155]), .B(_7725_), .Y(_7726_) );
	INVX1 INVX1_1001 ( .A(wSelec[158]), .Y(_7727_) );
	NAND2X1 NAND2X1_1615 ( .A(wSelec[157]), .B(_7727_), .Y(_7728_) );
	NOR2X1 NOR2X1_925 ( .A(_7726_), .B(_7728_), .Y(_7729_) );
	NOR2X1 NOR2X1_926 ( .A(wSelec[156]), .B(wSelec[155]), .Y(_7730_) );
	INVX1 INVX1_1002 ( .A(_7730_), .Y(_7731_) );
	NOR2X1 NOR2X1_927 ( .A(_7728_), .B(_7731_), .Y(_7732_) );
	AOI22X1 AOI22X1_1237 ( .A(wData[20]), .B(_7729_), .C(_7732_), .D(wData[16]), .Y(_7733_) );
	INVX1 INVX1_1003 ( .A(wSelec[155]), .Y(_7734_) );
	NAND2X1 NAND2X1_1616 ( .A(wSelec[156]), .B(_7734_), .Y(_7735_) );
	NOR2X1 NOR2X1_928 ( .A(_7735_), .B(_7728_), .Y(_7736_) );
	NAND2X1 NAND2X1_1617 ( .A(wData[24]), .B(_7736_), .Y(_7737_) );
	INVX1 INVX1_1004 ( .A(wSelec[157]), .Y(_7738_) );
	NAND2X1 NAND2X1_1618 ( .A(_7738_), .B(_7727_), .Y(_7739_) );
	NOR2X1 NOR2X1_929 ( .A(_7726_), .B(_7739_), .Y(_7740_) );
	NAND2X1 NAND2X1_1619 ( .A(wSelec[156]), .B(wSelec[155]), .Y(_7741_) );
	NOR2X1 NOR2X1_930 ( .A(_7741_), .B(_7728_), .Y(_7742_) );
	AOI22X1 AOI22X1_1238 ( .A(_7742_), .B(wData[28]), .C(wData[4]), .D(_7740_), .Y(_7743_) );
	NAND3X1 NAND3X1_383 ( .A(_7737_), .B(_7743_), .C(_7733_), .Y(_7744_) );
	NAND2X1 NAND2X1_1620 ( .A(wSelec[158]), .B(_7738_), .Y(_7745_) );
	NOR2X1 NOR2X1_931 ( .A(_7745_), .B(_7731_), .Y(_7746_) );
	NAND2X1 NAND2X1_1621 ( .A(wData[32]), .B(_7746_), .Y(_7747_) );
	NAND2X1 NAND2X1_1622 ( .A(wSelec[157]), .B(wSelec[158]), .Y(_7748_) );
	NOR2X1 NOR2X1_932 ( .A(_7748_), .B(_7735_), .Y(_7749_) );
	NOR2X1 NOR2X1_933 ( .A(_7748_), .B(_7726_), .Y(_7750_) );
	AOI22X1 AOI22X1_1239 ( .A(_7749_), .B(wData[56]), .C(wData[52]), .D(_7750_), .Y(_7751_) );
	NOR2X1 NOR2X1_934 ( .A(_7741_), .B(_7748_), .Y(_7752_) );
	NOR2X1 NOR2X1_935 ( .A(_7741_), .B(_7745_), .Y(_7753_) );
	AOI22X1 AOI22X1_1240 ( .A(wData[60]), .B(_7752_), .C(_7753_), .D(wData[44]), .Y(_7754_) );
	NAND3X1 NAND3X1_384 ( .A(_7747_), .B(_7754_), .C(_7751_), .Y(_7755_) );
	NOR2X1 NOR2X1_936 ( .A(_7735_), .B(_7745_), .Y(_7756_) );
	NAND2X1 NAND2X1_1623 ( .A(wData[40]), .B(_7756_), .Y(_7757_) );
	NOR2X1 NOR2X1_937 ( .A(_7745_), .B(_7726_), .Y(_7758_) );
	NAND2X1 NAND2X1_1624 ( .A(wData[36]), .B(_7758_), .Y(_7759_) );
	NOR2X1 NOR2X1_938 ( .A(_7739_), .B(_7731_), .Y(_7760_) );
	NAND2X1 NAND2X1_1625 ( .A(wData[0]), .B(_7760_), .Y(_7761_) );
	NAND3X1 NAND3X1_385 ( .A(_7757_), .B(_7759_), .C(_7761_), .Y(_7762_) );
	INVX1 INVX1_1005 ( .A(wData[48]), .Y(_7763_) );
	NOR2X1 NOR2X1_939 ( .A(_7738_), .B(_7727_), .Y(_7764_) );
	NAND2X1 NAND2X1_1626 ( .A(_7730_), .B(_7764_), .Y(_7765_) );
	NOR2X1 NOR2X1_940 ( .A(_7735_), .B(_7739_), .Y(_7766_) );
	NOR2X1 NOR2X1_941 ( .A(_7741_), .B(_7739_), .Y(_7767_) );
	AOI22X1 AOI22X1_1241 ( .A(_7766_), .B(wData[8]), .C(wData[12]), .D(_7767_), .Y(_7768_) );
	OAI21X1 OAI21X1_263 ( .A(_7763_), .B(_7765_), .C(_7768_), .Y(_7769_) );
	OR2X2 OR2X2_91 ( .A(_7769_), .B(_7762_), .Y(_7770_) );
	NOR3X1 NOR3X1_681 ( .A(_7744_), .B(_7755_), .C(_7770_), .Y(_7771_) );
	AND2X2 AND2X2_172 ( .A(_7771_), .B(_7535_), .Y(_7772_) );
	AOI21X1 AOI21X1_186 ( .A(_7626_), .B(_7724_), .C(_7772_), .Y(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_0_) );
	INVX1 INVX1_1006 ( .A(_7643_), .Y(_7773_) );
	AOI21X1 AOI21X1_187 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_7773_), .C(_7535_), .Y(_7774_) );
	AOI22X1 AOI22X1_1242 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_7543_), .C(_7559_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_7775_) );
	AOI22X1 AOI22X1_1243 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_7563_), .C(_7569_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_7776_) );
	NAND3X1 NAND3X1_386 ( .A(_7774_), .B(_7775_), .C(_7776_), .Y(_7777_) );
	INVX1 INVX1_1007 ( .A(_7603_), .Y(_7778_) );
	AOI22X1 AOI22X1_1244 ( .A(_7628_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_7778_), .Y(_7779_) );
	AOI22X1 AOI22X1_1245 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_7702_), .C(_7581_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_7780_) );
	INVX1 INVX1_1008 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_7781_) );
	INVX1 INVX1_1009 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_7782_) );
	OAI22X1 OAI22X1_213 ( .A(_7781_), .B(_7590_), .C(_7588_), .D(_7782_), .Y(_7783_) );
	INVX1 INVX1_1010 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_7784_) );
	NAND2X1 NAND2X1_1627 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_7691_), .Y(_7785_) );
	OAI21X1 OAI21X1_264 ( .A(_7784_), .B(_7596_), .C(_7785_), .Y(_7786_) );
	NOR2X1 NOR2X1_942 ( .A(_7783_), .B(_7786_), .Y(_7787_) );
	NAND3X1 NAND3X1_387 ( .A(_7779_), .B(_7780_), .C(_7787_), .Y(_7788_) );
	INVX1 INVX1_1011 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_7789_) );
	NAND2X1 NAND2X1_1628 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_7575_), .Y(_7790_) );
	OAI21X1 OAI21X1_265 ( .A(_7789_), .B(_7605_), .C(_7790_), .Y(_7791_) );
	INVX1 INVX1_1012 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_7792_) );
	INVX1 INVX1_1013 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_7793_) );
	OAI22X1 OAI22X1_214 ( .A(_7792_), .B(_7611_), .C(_7609_), .D(_7793_), .Y(_7794_) );
	NOR2X1 NOR2X1_943 ( .A(_7794_), .B(_7791_), .Y(_7795_) );
	AOI22X1 AOI22X1_1246 ( .A(_7695_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_7668_), .Y(_7796_) );
	AND2X2 AND2X2_173 ( .A(_7542_), .B(_7557_), .Y(_7797_) );
	AOI22X1 AOI22X1_1247 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_7667_), .C(_7797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_7798_) );
	NAND3X1 NAND3X1_388 ( .A(_7796_), .B(_7798_), .C(_7795_), .Y(_7799_) );
	NOR3X1 NOR3X1_682 ( .A(_7799_), .B(_7777_), .C(_7788_), .Y(_7800_) );
	INVX1 INVX1_1014 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_7801_) );
	NAND2X1 NAND2X1_1629 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_7630_), .Y(_7802_) );
	OAI21X1 OAI21X1_266 ( .A(_7632_), .B(_7801_), .C(_7802_), .Y(_7803_) );
	AOI21X1 AOI21X1_188 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_7679_), .C(_7803_), .Y(_7804_) );
	INVX1 INVX1_1015 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_7805_) );
	INVX1 INVX1_1016 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_7806_) );
	OAI22X1 OAI22X1_215 ( .A(_7806_), .B(_7638_), .C(_7639_), .D(_7805_), .Y(_7807_) );
	INVX1 INVX1_1017 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_7808_) );
	NAND2X1 NAND2X1_1630 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_7648_), .Y(_7809_) );
	OAI21X1 OAI21X1_267 ( .A(_7549_), .B(_7808_), .C(_7809_), .Y(_7810_) );
	NOR2X1 NOR2X1_944 ( .A(_7810_), .B(_7807_), .Y(_7811_) );
	INVX1 INVX1_1018 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_7812_) );
	INVX1 INVX1_1019 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_7813_) );
	OAI22X1 OAI22X1_216 ( .A(_7644_), .B(_7813_), .C(_7650_), .D(_7812_), .Y(_7814_) );
	INVX1 INVX1_1020 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_7815_) );
	NOR2X1 NOR2X1_945 ( .A(_7815_), .B(_7655_), .Y(_7816_) );
	INVX1 INVX1_1021 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_7817_) );
	NOR2X1 NOR2X1_946 ( .A(_7817_), .B(_7656_), .Y(_7818_) );
	NOR3X1 NOR3X1_683 ( .A(_7816_), .B(_7814_), .C(_7818_), .Y(_7819_) );
	NAND3X1 NAND3X1_389 ( .A(_7811_), .B(_7804_), .C(_7819_), .Y(_7820_) );
	AOI22X1 AOI22X1_1248 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_7660_), .C(_7661_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_7821_) );
	AOI22X1 AOI22X1_1249 ( .A(_7663_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_7664_), .Y(_7822_) );
	NAND2X1 NAND2X1_1631 ( .A(_7821_), .B(_7822_), .Y(_7823_) );
	AOI22X1 AOI22X1_1250 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_7671_), .C(_7670_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_7824_) );
	AOI22X1 AOI22X1_1251 ( .A(_7614_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_7621_), .Y(_7825_) );
	NAND2X1 NAND2X1_1632 ( .A(_7824_), .B(_7825_), .Y(_7826_) );
	NOR2X1 NOR2X1_947 ( .A(_7823_), .B(_7826_), .Y(_7827_) );
	AOI22X1 AOI22X1_1252 ( .A(_7675_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_7676_), .Y(_7828_) );
	AOI22X1 AOI22X1_1253 ( .A(_7577_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_7678_), .Y(_7829_) );
	NAND2X1 NAND2X1_1633 ( .A(_7828_), .B(_7829_), .Y(_7830_) );
	AOI22X1 AOI22X1_1254 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_7682_), .C(_7683_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_7831_) );
	AOI22X1 AOI22X1_1255 ( .A(_7685_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_7686_), .Y(_7832_) );
	NAND2X1 NAND2X1_1634 ( .A(_7832_), .B(_7831_), .Y(_7833_) );
	NOR2X1 NOR2X1_948 ( .A(_7830_), .B(_7833_), .Y(_7834_) );
	NAND2X1 NAND2X1_1635 ( .A(_7834_), .B(_7827_), .Y(_7835_) );
	AOI22X1 AOI22X1_1256 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_7692_), .C(_7593_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_7836_) );
	AOI22X1 AOI22X1_1257 ( .A(_7616_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_7694_), .Y(_7837_) );
	NAND2X1 NAND2X1_1636 ( .A(_7836_), .B(_7837_), .Y(_7838_) );
	AOI22X1 AOI22X1_1258 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_7583_), .C(_7703_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_7839_) );
	NAND2X1 NAND2X1_1637 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_7698_), .Y(_7840_) );
	NAND2X1 NAND2X1_1638 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_7700_), .Y(_7841_) );
	NAND3X1 NAND3X1_390 ( .A(_7840_), .B(_7841_), .C(_7839_), .Y(_7842_) );
	NOR2X1 NOR2X1_949 ( .A(_7842_), .B(_7838_), .Y(_7843_) );
	AOI22X1 AOI22X1_1259 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_7707_), .C(_7708_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_7844_) );
	NAND2X1 NAND2X1_1639 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_7710_), .Y(_7845_) );
	NAND2X1 NAND2X1_1640 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_7712_), .Y(_7846_) );
	NAND3X1 NAND3X1_391 ( .A(_7845_), .B(_7846_), .C(_7844_), .Y(_7847_) );
	AOI22X1 AOI22X1_1260 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_7716_), .C(_7715_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_7848_) );
	AOI22X1 AOI22X1_1261 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_7719_), .C(_7718_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_7849_) );
	NAND2X1 NAND2X1_1641 ( .A(_7848_), .B(_7849_), .Y(_7850_) );
	NOR2X1 NOR2X1_950 ( .A(_7850_), .B(_7847_), .Y(_7851_) );
	NAND2X1 NAND2X1_1642 ( .A(_7843_), .B(_7851_), .Y(_7852_) );
	NOR3X1 NOR3X1_684 ( .A(_7835_), .B(_7820_), .C(_7852_), .Y(_7853_) );
	AOI21X1 AOI21X1_189 ( .A(wData[21]), .B(_7729_), .C(_7534_), .Y(_7854_) );
	AOI22X1 AOI22X1_1262 ( .A(_7732_), .B(wData[17]), .C(wData[1]), .D(_7760_), .Y(_7855_) );
	AOI22X1 AOI22X1_1263 ( .A(_7753_), .B(wData[45]), .C(wData[25]), .D(_7736_), .Y(_7856_) );
	NAND3X1 NAND3X1_392 ( .A(_7854_), .B(_7856_), .C(_7855_), .Y(_7857_) );
	NAND3X1 NAND3X1_393 ( .A(wData[49]), .B(_7730_), .C(_7764_), .Y(_7858_) );
	AOI22X1 AOI22X1_1264 ( .A(wData[61]), .B(_7752_), .C(_7740_), .D(wData[5]), .Y(_7859_) );
	AND2X2 AND2X2_174 ( .A(_7859_), .B(_7858_), .Y(_7860_) );
	AOI22X1 AOI22X1_1265 ( .A(_7749_), .B(wData[57]), .C(wData[41]), .D(_7756_), .Y(_7861_) );
	AOI22X1 AOI22X1_1266 ( .A(wData[53]), .B(_7750_), .C(_7746_), .D(wData[33]), .Y(_7862_) );
	AND2X2 AND2X2_175 ( .A(_7862_), .B(_7861_), .Y(_7863_) );
	AOI22X1 AOI22X1_1267 ( .A(_7766_), .B(wData[9]), .C(wData[13]), .D(_7767_), .Y(_7864_) );
	AOI22X1 AOI22X1_1268 ( .A(_7742_), .B(wData[29]), .C(wData[37]), .D(_7758_), .Y(_7865_) );
	AND2X2 AND2X2_176 ( .A(_7864_), .B(_7865_), .Y(_7866_) );
	NAND3X1 NAND3X1_394 ( .A(_7860_), .B(_7866_), .C(_7863_), .Y(_7867_) );
	NOR2X1 NOR2X1_951 ( .A(_7857_), .B(_7867_), .Y(_7868_) );
	AOI21X1 AOI21X1_190 ( .A(_7800_), .B(_7853_), .C(_7868_), .Y(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_1_) );
	AOI21X1 AOI21X1_191 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_7773_), .C(_7535_), .Y(_7869_) );
	INVX1 INVX1_1022 ( .A(_7632_), .Y(_7870_) );
	AOI22X1 AOI22X1_1269 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_7543_), .C(_7870_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_7871_) );
	INVX1 INVX1_1023 ( .A(_7644_), .Y(_7872_) );
	AOI22X1 AOI22X1_1270 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_7679_), .C(_7872_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_7873_) );
	NAND3X1 NAND3X1_395 ( .A(_7873_), .B(_7869_), .C(_7871_), .Y(_7874_) );
	AOI22X1 AOI22X1_1271 ( .A(_7628_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_7778_), .Y(_7875_) );
	AOI22X1 AOI22X1_1272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_7577_), .C(_7550_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_7876_) );
	INVX1 INVX1_1024 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_7877_) );
	NAND2X1 NAND2X1_1643 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_7667_), .Y(_7878_) );
	OAI21X1 OAI21X1_268 ( .A(_7877_), .B(_7639_), .C(_7878_), .Y(_7879_) );
	INVX1 INVX1_1025 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_7880_) );
	NAND2X1 NAND2X1_1644 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_7593_), .Y(_7881_) );
	OAI21X1 OAI21X1_269 ( .A(_7880_), .B(_7596_), .C(_7881_), .Y(_7882_) );
	NOR2X1 NOR2X1_952 ( .A(_7879_), .B(_7882_), .Y(_7883_) );
	NAND3X1 NAND3X1_396 ( .A(_7875_), .B(_7876_), .C(_7883_), .Y(_7884_) );
	INVX1 INVX1_1026 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_7885_) );
	NAND2X1 NAND2X1_1645 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_7575_), .Y(_7886_) );
	OAI21X1 OAI21X1_270 ( .A(_7885_), .B(_7605_), .C(_7886_), .Y(_7887_) );
	INVX1 INVX1_1027 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_7888_) );
	INVX1 INVX1_1028 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_7889_) );
	OAI22X1 OAI22X1_217 ( .A(_7888_), .B(_7611_), .C(_7609_), .D(_7889_), .Y(_7890_) );
	NOR2X1 NOR2X1_953 ( .A(_7890_), .B(_7887_), .Y(_7891_) );
	AOI22X1 AOI22X1_1273 ( .A(_7695_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_7668_), .Y(_7892_) );
	AND2X2 AND2X2_177 ( .A(_7567_), .B(_7589_), .Y(_7893_) );
	AOI22X1 AOI22X1_1274 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_7893_), .C(_7797_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_7894_) );
	NAND3X1 NAND3X1_397 ( .A(_7892_), .B(_7894_), .C(_7891_), .Y(_7895_) );
	NOR3X1 NOR3X1_685 ( .A(_7895_), .B(_7874_), .C(_7884_), .Y(_7896_) );
	INVX1 INVX1_1029 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_7897_) );
	NOR3X1 NOR3X1_686 ( .A(_7897_), .B(_7562_), .C(_7561_), .Y(_7898_) );
	AND2X2 AND2X2_178 ( .A(_7583_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_7899_) );
	AND2X2 AND2X2_179 ( .A(_7703_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_7900_) );
	NOR3X1 NOR3X1_687 ( .A(_7900_), .B(_7899_), .C(_7898_), .Y(_7901_) );
	INVX1 INVX1_1030 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_7902_) );
	INVX1 INVX1_1031 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_7903_) );
	OAI22X1 OAI22X1_218 ( .A(_7903_), .B(_7638_), .C(_7588_), .D(_7902_), .Y(_7904_) );
	INVX1 INVX1_1032 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_7905_) );
	INVX1 INVX1_1033 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_7906_) );
	NAND2X1 NAND2X1_1646 ( .A(_7579_), .B(_7580_), .Y(_7907_) );
	OAI22X1 OAI22X1_219 ( .A(_7907_), .B(_7906_), .C(_7905_), .D(_7558_), .Y(_7908_) );
	NOR2X1 NOR2X1_954 ( .A(_7904_), .B(_7908_), .Y(_7909_) );
	INVX1 INVX1_1034 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_7910_) );
	NOR3X1 NOR3X1_688 ( .A(_7539_), .B(_7556_), .C(_7547_), .Y(_7911_) );
	NAND2X1 NAND2X1_1647 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_7911_), .Y(_7912_) );
	OAI21X1 OAI21X1_271 ( .A(_7568_), .B(_7910_), .C(_7912_), .Y(_7913_) );
	INVX1 INVX1_1035 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_7914_) );
	INVX1 INVX1_1036 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_7915_) );
	OAI22X1 OAI22X1_220 ( .A(_7655_), .B(_7915_), .C(_7914_), .D(_7656_), .Y(_7916_) );
	NOR2X1 NOR2X1_955 ( .A(_7913_), .B(_7916_), .Y(_7917_) );
	NAND3X1 NAND3X1_398 ( .A(_7901_), .B(_7917_), .C(_7909_), .Y(_7918_) );
	AOI22X1 AOI22X1_1275 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_7660_), .C(_7661_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_7919_) );
	AOI22X1 AOI22X1_1276 ( .A(_7663_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_7664_), .Y(_7920_) );
	NAND2X1 NAND2X1_1648 ( .A(_7919_), .B(_7920_), .Y(_7921_) );
	AOI22X1 AOI22X1_1277 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_7671_), .C(_7670_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_7922_) );
	AOI22X1 AOI22X1_1278 ( .A(_7614_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_7621_), .Y(_7923_) );
	NAND2X1 NAND2X1_1649 ( .A(_7922_), .B(_7923_), .Y(_7924_) );
	NOR2X1 NOR2X1_956 ( .A(_7921_), .B(_7924_), .Y(_7925_) );
	AOI22X1 AOI22X1_1279 ( .A(_7675_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_7676_), .Y(_7926_) );
	AOI22X1 AOI22X1_1280 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_7702_), .C(_7678_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_7927_) );
	NAND2X1 NAND2X1_1650 ( .A(_7927_), .B(_7926_), .Y(_7928_) );
	AOI22X1 AOI22X1_1281 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_7682_), .C(_7683_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_7929_) );
	AOI22X1 AOI22X1_1282 ( .A(_7685_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_7686_), .Y(_7930_) );
	NAND2X1 NAND2X1_1651 ( .A(_7930_), .B(_7929_), .Y(_7931_) );
	NOR2X1 NOR2X1_957 ( .A(_7928_), .B(_7931_), .Y(_7932_) );
	NAND2X1 NAND2X1_1652 ( .A(_7932_), .B(_7925_), .Y(_7933_) );
	AOI22X1 AOI22X1_1283 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_7692_), .C(_7691_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_7934_) );
	AOI22X1 AOI22X1_1284 ( .A(_7616_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_7694_), .Y(_7935_) );
	NAND2X1 NAND2X1_1653 ( .A(_7934_), .B(_7935_), .Y(_7936_) );
	AOI22X1 AOI22X1_1285 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_7700_), .C(_7698_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_7937_) );
	AOI22X1 AOI22X1_1286 ( .A(_7630_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_7648_), .Y(_7938_) );
	NAND2X1 NAND2X1_1654 ( .A(_7938_), .B(_7937_), .Y(_7939_) );
	NOR2X1 NOR2X1_958 ( .A(_7939_), .B(_7936_), .Y(_7940_) );
	AOI22X1 AOI22X1_1287 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_7707_), .C(_7708_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_7941_) );
	NAND2X1 NAND2X1_1655 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_7710_), .Y(_7942_) );
	NAND2X1 NAND2X1_1656 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_7712_), .Y(_7943_) );
	NAND3X1 NAND3X1_399 ( .A(_7942_), .B(_7943_), .C(_7941_), .Y(_7944_) );
	AOI22X1 AOI22X1_1288 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_7716_), .C(_7715_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_7945_) );
	AOI22X1 AOI22X1_1289 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_7719_), .C(_7718_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_7946_) );
	NAND2X1 NAND2X1_1657 ( .A(_7945_), .B(_7946_), .Y(_7947_) );
	NOR2X1 NOR2X1_959 ( .A(_7947_), .B(_7944_), .Y(_7948_) );
	NAND2X1 NAND2X1_1658 ( .A(_7940_), .B(_7948_), .Y(_7949_) );
	NOR3X1 NOR3X1_689 ( .A(_7933_), .B(_7918_), .C(_7949_), .Y(_7950_) );
	AOI22X1 AOI22X1_1290 ( .A(_7756_), .B(wData[42]), .C(wData[38]), .D(_7758_), .Y(_7951_) );
	AOI22X1 AOI22X1_1291 ( .A(_7753_), .B(wData[46]), .C(_7760_), .D(wData[2]), .Y(_7952_) );
	NAND2X1 NAND2X1_1659 ( .A(_7951_), .B(_7952_), .Y(_7953_) );
	AOI21X1 AOI21X1_192 ( .A(wData[34]), .B(_7746_), .C(_7953_), .Y(_7954_) );
	INVX1 INVX1_1037 ( .A(wData[50]), .Y(_7955_) );
	AOI22X1 AOI22X1_1292 ( .A(_7766_), .B(wData[10]), .C(wData[14]), .D(_7767_), .Y(_7956_) );
	OAI21X1 OAI21X1_272 ( .A(_7955_), .B(_7765_), .C(_7956_), .Y(_7957_) );
	AOI22X1 AOI22X1_1293 ( .A(_7729_), .B(wData[22]), .C(wData[18]), .D(_7732_), .Y(_7958_) );
	NAND2X1 NAND2X1_1660 ( .A(wData[26]), .B(_7736_), .Y(_7959_) );
	AOI22X1 AOI22X1_1294 ( .A(_7742_), .B(wData[30]), .C(wData[6]), .D(_7740_), .Y(_7960_) );
	NAND3X1 NAND3X1_400 ( .A(_7959_), .B(_7960_), .C(_7958_), .Y(_7961_) );
	NOR2X1 NOR2X1_960 ( .A(_7957_), .B(_7961_), .Y(_7962_) );
	NAND2X1 NAND2X1_1661 ( .A(wData[58]), .B(_7749_), .Y(_7963_) );
	NAND2X1 NAND2X1_1662 ( .A(wData[54]), .B(_7750_), .Y(_7964_) );
	NAND2X1 NAND2X1_1663 ( .A(_7963_), .B(_7964_), .Y(_7965_) );
	AOI21X1 AOI21X1_193 ( .A(wData[62]), .B(_7752_), .C(_7965_), .Y(_7966_) );
	NAND3X1 NAND3X1_401 ( .A(_7954_), .B(_7966_), .C(_7962_), .Y(_7967_) );
	NOR2X1 NOR2X1_961 ( .A(_7534_), .B(_7967_), .Y(_7968_) );
	AOI21X1 AOI21X1_194 ( .A(_7896_), .B(_7950_), .C(_7968_), .Y(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_2_) );
	AOI21X1 AOI21X1_195 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_7778_), .C(_7535_), .Y(_7969_) );
	AOI22X1 AOI22X1_1295 ( .A(_7550_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_7870_), .Y(_7970_) );
	AOI22X1 AOI22X1_1296 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_7872_), .C(_7628_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_7971_) );
	NAND3X1 NAND3X1_402 ( .A(_7971_), .B(_7969_), .C(_7970_), .Y(_7972_) );
	AOI22X1 AOI22X1_1297 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_7577_), .C(_7575_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_7973_) );
	AOI22X1 AOI22X1_1298 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_7648_), .C(_7773_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_7974_) );
	INVX1 INVX1_1038 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_7975_) );
	INVX1 INVX1_1039 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_7976_) );
	OAI22X1 OAI22X1_221 ( .A(_7975_), .B(_7590_), .C(_7639_), .D(_7976_), .Y(_7977_) );
	INVX1 INVX1_1040 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_7978_) );
	NAND2X1 NAND2X1_1664 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_7691_), .Y(_7979_) );
	OAI21X1 OAI21X1_273 ( .A(_7978_), .B(_7596_), .C(_7979_), .Y(_7980_) );
	NOR2X1 NOR2X1_962 ( .A(_7977_), .B(_7980_), .Y(_7981_) );
	NAND3X1 NAND3X1_403 ( .A(_7973_), .B(_7974_), .C(_7981_), .Y(_7982_) );
	AND2X2 AND2X2_180 ( .A(_7604_), .B(_7538_), .Y(_7983_) );
	AOI22X1 AOI22X1_1299 ( .A(_7543_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_7983_), .Y(_7984_) );
	AND2X2 AND2X2_181 ( .A(_7602_), .B(_7567_), .Y(_7985_) );
	AND2X2 AND2X2_182 ( .A(_7610_), .B(_7567_), .Y(_7986_) );
	AOI22X1 AOI22X1_1300 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_7986_), .C(_7985_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_7987_) );
	NAND2X1 NAND2X1_1665 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_7695_), .Y(_7988_) );
	NAND2X1 NAND2X1_1666 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_7668_), .Y(_7989_) );
	NAND2X1 NAND2X1_1667 ( .A(_7988_), .B(_7989_), .Y(_7990_) );
	INVX1 INVX1_1041 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_7991_) );
	NAND2X1 NAND2X1_1668 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_7667_), .Y(_7992_) );
	OAI21X1 OAI21X1_274 ( .A(_7991_), .B(_7620_), .C(_7992_), .Y(_7993_) );
	NOR2X1 NOR2X1_963 ( .A(_7990_), .B(_7993_), .Y(_7994_) );
	NAND3X1 NAND3X1_404 ( .A(_7984_), .B(_7987_), .C(_7994_), .Y(_7995_) );
	NOR3X1 NOR3X1_690 ( .A(_7982_), .B(_7972_), .C(_7995_), .Y(_7996_) );
	INVX1 INVX1_1042 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_7997_) );
	NAND2X1 NAND2X1_1669 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_7583_), .Y(_7998_) );
	OAI21X1 OAI21X1_275 ( .A(_7588_), .B(_7997_), .C(_7998_), .Y(_7999_) );
	AOI21X1 AOI21X1_196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_7563_), .C(_7999_), .Y(_8000_) );
	INVX1 INVX1_1043 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_8001_) );
	INVX1 INVX1_1044 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_8002_) );
	OAI22X1 OAI22X1_222 ( .A(_7907_), .B(_8002_), .C(_8001_), .D(_7558_), .Y(_8003_) );
	INVX1 INVX1_1045 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_8004_) );
	NAND2X1 NAND2X1_1670 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_7703_), .Y(_8005_) );
	OAI21X1 OAI21X1_276 ( .A(_7568_), .B(_8004_), .C(_8005_), .Y(_8006_) );
	NOR2X1 NOR2X1_964 ( .A(_8006_), .B(_8003_), .Y(_8007_) );
	INVX1 INVX1_1046 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_8008_) );
	INVX1 INVX1_1047 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_8009_) );
	OAI22X1 OAI22X1_223 ( .A(_7655_), .B(_8009_), .C(_8008_), .D(_7656_), .Y(_8010_) );
	INVX1 INVX1_1048 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_8011_) );
	NAND2X1 NAND2X1_1671 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_7702_), .Y(_8012_) );
	OAI21X1 OAI21X1_277 ( .A(_8011_), .B(_7638_), .C(_8012_), .Y(_8013_) );
	NOR2X1 NOR2X1_965 ( .A(_8013_), .B(_8010_), .Y(_8014_) );
	NAND3X1 NAND3X1_405 ( .A(_8000_), .B(_8014_), .C(_8007_), .Y(_8015_) );
	AOI22X1 AOI22X1_1301 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_7660_), .C(_7661_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_8016_) );
	AOI22X1 AOI22X1_1302 ( .A(_7663_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_7664_), .Y(_8017_) );
	NAND2X1 NAND2X1_1672 ( .A(_8016_), .B(_8017_), .Y(_8018_) );
	AOI22X1 AOI22X1_1303 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_7671_), .C(_7670_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_8019_) );
	AOI22X1 AOI22X1_1304 ( .A(_7614_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_7621_), .Y(_8020_) );
	NAND2X1 NAND2X1_1673 ( .A(_8019_), .B(_8020_), .Y(_8021_) );
	NOR2X1 NOR2X1_966 ( .A(_8018_), .B(_8021_), .Y(_8022_) );
	AOI22X1 AOI22X1_1305 ( .A(_7675_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_7676_), .Y(_8023_) );
	AOI22X1 AOI22X1_1306 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_7911_), .C(_7678_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_8024_) );
	NAND2X1 NAND2X1_1674 ( .A(_8024_), .B(_8023_), .Y(_8025_) );
	AOI22X1 AOI22X1_1307 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_7682_), .C(_7683_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_8026_) );
	AOI22X1 AOI22X1_1308 ( .A(_7685_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_7686_), .Y(_8027_) );
	NAND2X1 NAND2X1_1675 ( .A(_8027_), .B(_8026_), .Y(_8028_) );
	NOR2X1 NOR2X1_967 ( .A(_8025_), .B(_8028_), .Y(_8029_) );
	NAND2X1 NAND2X1_1676 ( .A(_8029_), .B(_8022_), .Y(_8030_) );
	AOI22X1 AOI22X1_1309 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_7692_), .C(_7593_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_8031_) );
	AOI22X1 AOI22X1_1310 ( .A(_7616_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_7694_), .Y(_8032_) );
	NAND2X1 NAND2X1_1677 ( .A(_8031_), .B(_8032_), .Y(_8033_) );
	AOI22X1 AOI22X1_1311 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_7700_), .C(_7698_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_8034_) );
	AOI22X1 AOI22X1_1312 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_7630_), .C(_7679_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_8035_) );
	NAND2X1 NAND2X1_1678 ( .A(_8035_), .B(_8034_), .Y(_8036_) );
	NOR2X1 NOR2X1_968 ( .A(_8036_), .B(_8033_), .Y(_8037_) );
	AOI22X1 AOI22X1_1313 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_7707_), .C(_7708_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_8038_) );
	NAND2X1 NAND2X1_1679 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_7710_), .Y(_8039_) );
	NAND2X1 NAND2X1_1680 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_7712_), .Y(_8040_) );
	NAND3X1 NAND3X1_406 ( .A(_8039_), .B(_8040_), .C(_8038_), .Y(_8041_) );
	AOI22X1 AOI22X1_1314 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_7716_), .C(_7715_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_8042_) );
	AOI22X1 AOI22X1_1315 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_7719_), .C(_7718_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_8043_) );
	NAND2X1 NAND2X1_1681 ( .A(_8042_), .B(_8043_), .Y(_8044_) );
	NOR2X1 NOR2X1_969 ( .A(_8044_), .B(_8041_), .Y(_8045_) );
	NAND2X1 NAND2X1_1682 ( .A(_8037_), .B(_8045_), .Y(_8046_) );
	NOR3X1 NOR3X1_691 ( .A(_8030_), .B(_8015_), .C(_8046_), .Y(_8047_) );
	NAND2X1 NAND2X1_1683 ( .A(wData[59]), .B(_7749_), .Y(_8048_) );
	OAI21X1 OAI21X1_278 ( .A(_7533_), .B(wBusy_bF_buf3), .C(_8048_), .Y(_8049_) );
	NAND2X1 NAND2X1_1684 ( .A(wData[7]), .B(_7740_), .Y(_8050_) );
	NAND2X1 NAND2X1_1685 ( .A(wData[55]), .B(_7750_), .Y(_8051_) );
	AOI22X1 AOI22X1_1316 ( .A(wData[63]), .B(_7752_), .C(_7742_), .D(wData[31]), .Y(_8052_) );
	NAND3X1 NAND3X1_407 ( .A(_8050_), .B(_8051_), .C(_8052_), .Y(_8053_) );
	OR2X2 OR2X2_92 ( .A(_8053_), .B(_8049_), .Y(_8054_) );
	INVX1 INVX1_1049 ( .A(wData[51]), .Y(_8055_) );
	NAND2X1 NAND2X1_1686 ( .A(wData[47]), .B(_7753_), .Y(_8056_) );
	OAI21X1 OAI21X1_279 ( .A(_8055_), .B(_7765_), .C(_8056_), .Y(_8057_) );
	AOI21X1 AOI21X1_197 ( .A(wData[3]), .B(_7760_), .C(_8057_), .Y(_8058_) );
	AOI22X1 AOI22X1_1317 ( .A(_7766_), .B(wData[11]), .C(wData[15]), .D(_7767_), .Y(_8059_) );
	AOI22X1 AOI22X1_1318 ( .A(_7729_), .B(wData[23]), .C(wData[27]), .D(_7736_), .Y(_8060_) );
	AND2X2 AND2X2_183 ( .A(_8059_), .B(_8060_), .Y(_8061_) );
	NAND2X1 NAND2X1_1687 ( .A(wData[39]), .B(_7758_), .Y(_8062_) );
	NAND2X1 NAND2X1_1688 ( .A(wData[43]), .B(_7756_), .Y(_8063_) );
	NAND2X1 NAND2X1_1689 ( .A(_8062_), .B(_8063_), .Y(_8064_) );
	NAND2X1 NAND2X1_1690 ( .A(wData[19]), .B(_7732_), .Y(_8065_) );
	NAND2X1 NAND2X1_1691 ( .A(wData[35]), .B(_7746_), .Y(_8066_) );
	NAND2X1 NAND2X1_1692 ( .A(_8065_), .B(_8066_), .Y(_8067_) );
	NOR2X1 NOR2X1_970 ( .A(_8064_), .B(_8067_), .Y(_8068_) );
	NAND3X1 NAND3X1_408 ( .A(_8061_), .B(_8058_), .C(_8068_), .Y(_8069_) );
	NOR2X1 NOR2X1_971 ( .A(_8054_), .B(_8069_), .Y(_8070_) );
	AOI21X1 AOI21X1_198 ( .A(_7996_), .B(_8047_), .C(_8070_), .Y(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_3_) );
	INVX1 INVX1_1050 ( .A(wSelec[165]), .Y(_8071_) );
	NOR2X1 NOR2X1_972 ( .A(wBusy_bF_buf2), .B(_8071_), .Y(_8072_) );
	INVX1 INVX1_1051 ( .A(_8072_), .Y(_8073_) );
	INVX1 INVX1_1052 ( .A(wSelec[175]), .Y(_8074_) );
	NAND2X1 NAND2X1_1693 ( .A(wSelec[174]), .B(_8074_), .Y(_8075_) );
	INVX2 INVX2_27 ( .A(_8075_), .Y(_8076_) );
	OR2X2 OR2X2_93 ( .A(wSelec[171]), .B(wSelec[170]), .Y(_8077_) );
	INVX1 INVX1_1053 ( .A(wSelec[173]), .Y(_8078_) );
	NAND2X1 NAND2X1_1694 ( .A(wSelec[172]), .B(_8078_), .Y(_8079_) );
	NOR2X1 NOR2X1_973 ( .A(_8077_), .B(_8079_), .Y(_8080_) );
	AND2X2 AND2X2_184 ( .A(_8080_), .B(_8076_), .Y(_8081_) );
	AOI21X1 AOI21X1_199 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_8081_), .C(_8073_), .Y(_8082_) );
	INVX1 INVX1_1054 ( .A(wSelec[171]), .Y(_8083_) );
	NAND2X1 NAND2X1_1695 ( .A(wSelec[170]), .B(_8083_), .Y(_8084_) );
	OR2X2 OR2X2_94 ( .A(wSelec[172]), .B(wSelec[173]), .Y(_8085_) );
	NOR2X1 NOR2X1_974 ( .A(_8085_), .B(_8084_), .Y(_8086_) );
	NAND2X1 NAND2X1_1696 ( .A(_8076_), .B(_8086_), .Y(_8087_) );
	INVX1 INVX1_1055 ( .A(_8087_), .Y(_8088_) );
	INVX1 INVX1_1056 ( .A(wSelec[170]), .Y(_8089_) );
	NAND2X1 NAND2X1_1697 ( .A(wSelec[171]), .B(_8089_), .Y(_8090_) );
	INVX1 INVX1_1057 ( .A(wSelec[172]), .Y(_8091_) );
	NAND2X1 NAND2X1_1698 ( .A(wSelec[173]), .B(_8091_), .Y(_8092_) );
	NOR2X1 NOR2X1_975 ( .A(_8090_), .B(_8092_), .Y(_8093_) );
	NAND2X1 NAND2X1_1699 ( .A(wSelec[174]), .B(wSelec[175]), .Y(_8094_) );
	INVX1 INVX1_1058 ( .A(_8094_), .Y(_8095_) );
	NAND2X1 NAND2X1_1700 ( .A(_8095_), .B(_8093_), .Y(_8096_) );
	INVX1 INVX1_1059 ( .A(_8096_), .Y(_8097_) );
	AOI22X1 AOI22X1_1319 ( .A(_8088_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_8097_), .Y(_8098_) );
	OR2X2 OR2X2_95 ( .A(_8084_), .B(_8085_), .Y(_8099_) );
	OR2X2 OR2X2_96 ( .A(wSelec[174]), .B(wSelec[175]), .Y(_8100_) );
	NOR2X1 NOR2X1_976 ( .A(_8100_), .B(_8099_), .Y(_8101_) );
	NOR2X1 NOR2X1_977 ( .A(_8079_), .B(_8084_), .Y(_8102_) );
	INVX1 INVX1_1060 ( .A(wSelec[174]), .Y(_8103_) );
	NAND2X1 NAND2X1_1701 ( .A(wSelec[175]), .B(_8103_), .Y(_8104_) );
	INVX2 INVX2_28 ( .A(_8104_), .Y(_8105_) );
	NAND2X1 NAND2X1_1702 ( .A(_8105_), .B(_8102_), .Y(_8106_) );
	INVX1 INVX1_1061 ( .A(_8106_), .Y(_8107_) );
	AOI22X1 AOI22X1_1320 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_8101_), .C(_8107_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_8108_) );
	NAND3X1 NAND3X1_409 ( .A(_8082_), .B(_8108_), .C(_8098_), .Y(_8109_) );
	NOR2X1 NOR2X1_978 ( .A(wSelec[171]), .B(wSelec[170]), .Y(_8110_) );
	NOR2X1 NOR2X1_979 ( .A(wSelec[172]), .B(wSelec[173]), .Y(_8111_) );
	NAND2X1 NAND2X1_1703 ( .A(_8110_), .B(_8111_), .Y(_8112_) );
	NOR2X1 NOR2X1_980 ( .A(_8075_), .B(_8112_), .Y(_8113_) );
	NAND2X1 NAND2X1_1704 ( .A(wSelec[171]), .B(wSelec[170]), .Y(_8114_) );
	NOR3X1 NOR3X1_692 ( .A(_8085_), .B(_8114_), .C(_8075_), .Y(_8115_) );
	AOI22X1 AOI22X1_1321 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_8115_), .C(_8113_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_8116_) );
	INVX1 INVX1_1062 ( .A(_8100_), .Y(_8117_) );
	NOR2X1 NOR2X1_981 ( .A(_8085_), .B(_8090_), .Y(_8118_) );
	AND2X2 AND2X2_185 ( .A(_8118_), .B(_8117_), .Y(_8119_) );
	NAND2X1 NAND2X1_1705 ( .A(wSelec[172]), .B(wSelec[173]), .Y(_8120_) );
	NOR3X1 NOR3X1_693 ( .A(_8094_), .B(_8114_), .C(_8120_), .Y(_8121_) );
	AOI22X1 AOI22X1_1322 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_8121_), .C(_8119_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_8122_) );
	INVX1 INVX1_1063 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_8123_) );
	INVX1 INVX1_1064 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_8124_) );
	NOR2X1 NOR2X1_982 ( .A(_8084_), .B(_8092_), .Y(_8125_) );
	NAND2X1 NAND2X1_1706 ( .A(_8095_), .B(_8125_), .Y(_8126_) );
	NOR2X1 NOR2X1_983 ( .A(_8114_), .B(_8120_), .Y(_8127_) );
	NAND2X1 NAND2X1_1707 ( .A(_8127_), .B(_8105_), .Y(_8128_) );
	OAI22X1 OAI22X1_224 ( .A(_8123_), .B(_8128_), .C(_8126_), .D(_8124_), .Y(_8129_) );
	INVX1 INVX1_1065 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_8130_) );
	NOR3X1 NOR3X1_694 ( .A(_8075_), .B(_8090_), .C(_8092_), .Y(_8131_) );
	NAND2X1 NAND2X1_1708 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_8131_), .Y(_8132_) );
	NOR2X1 NOR2X1_984 ( .A(_8114_), .B(_8079_), .Y(_8133_) );
	NAND2X1 NAND2X1_1709 ( .A(_8105_), .B(_8133_), .Y(_8134_) );
	OAI21X1 OAI21X1_280 ( .A(_8130_), .B(_8134_), .C(_8132_), .Y(_8135_) );
	NOR2X1 NOR2X1_985 ( .A(_8129_), .B(_8135_), .Y(_8136_) );
	NAND3X1 NAND3X1_410 ( .A(_8116_), .B(_8122_), .C(_8136_), .Y(_8137_) );
	INVX1 INVX1_1066 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_8138_) );
	INVX1 INVX1_1067 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_8139_) );
	NOR2X1 NOR2X1_986 ( .A(_8079_), .B(_8090_), .Y(_8140_) );
	NAND2X1 NAND2X1_1710 ( .A(_8076_), .B(_8140_), .Y(_8141_) );
	NOR2X1 NOR2X1_987 ( .A(_8077_), .B(_8092_), .Y(_8142_) );
	NAND2X1 NAND2X1_1711 ( .A(_8076_), .B(_8142_), .Y(_8143_) );
	OAI22X1 OAI22X1_225 ( .A(_8143_), .B(_8138_), .C(_8139_), .D(_8141_), .Y(_8144_) );
	INVX1 INVX1_1068 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_8145_) );
	INVX1 INVX1_1069 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_8146_) );
	NAND2X1 NAND2X1_1712 ( .A(_8105_), .B(_8140_), .Y(_8147_) );
	NOR2X1 NOR2X1_988 ( .A(_8114_), .B(_8085_), .Y(_8148_) );
	NAND2X1 NAND2X1_1713 ( .A(_8105_), .B(_8148_), .Y(_8149_) );
	OAI22X1 OAI22X1_226 ( .A(_8145_), .B(_8149_), .C(_8147_), .D(_8146_), .Y(_8150_) );
	NOR2X1 NOR2X1_989 ( .A(_8150_), .B(_8144_), .Y(_8151_) );
	NOR3X1 NOR3X1_695 ( .A(_8084_), .B(_8120_), .C(_8104_), .Y(_8152_) );
	NAND2X1 NAND2X1_1714 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_8152_), .Y(_8153_) );
	NOR3X1 NOR3X1_696 ( .A(_8092_), .B(_8114_), .C(_8104_), .Y(_8154_) );
	NAND2X1 NAND2X1_1715 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_8154_), .Y(_8155_) );
	NAND2X1 NAND2X1_1716 ( .A(_8153_), .B(_8155_), .Y(_8156_) );
	INVX1 INVX1_1070 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_8157_) );
	NAND2X1 NAND2X1_1717 ( .A(_8095_), .B(_8080_), .Y(_8158_) );
	NOR3X1 NOR3X1_697 ( .A(_8090_), .B(_8092_), .C(_8104_), .Y(_8159_) );
	NAND2X1 NAND2X1_1718 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_8159_), .Y(_8160_) );
	OAI21X1 OAI21X1_281 ( .A(_8157_), .B(_8158_), .C(_8160_), .Y(_8161_) );
	NOR2X1 NOR2X1_990 ( .A(_8156_), .B(_8161_), .Y(_8162_) );
	NAND2X1 NAND2X1_1719 ( .A(_8151_), .B(_8162_), .Y(_8163_) );
	NOR3X1 NOR3X1_698 ( .A(_8109_), .B(_8163_), .C(_8137_), .Y(_8164_) );
	NAND2X1 NAND2X1_1720 ( .A(_8076_), .B(_8133_), .Y(_8165_) );
	INVX1 INVX1_1071 ( .A(_8165_), .Y(_8166_) );
	INVX1 INVX1_1072 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_8167_) );
	NOR3X1 NOR3X1_699 ( .A(_8077_), .B(_8100_), .C(_8079_), .Y(_8168_) );
	NAND2X1 NAND2X1_1721 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_8168_), .Y(_8169_) );
	NAND2X1 NAND2X1_1722 ( .A(_8117_), .B(_8140_), .Y(_8170_) );
	OAI21X1 OAI21X1_282 ( .A(_8170_), .B(_8167_), .C(_8169_), .Y(_8171_) );
	AOI21X1 AOI21X1_200 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_8166_), .C(_8171_), .Y(_8172_) );
	INVX1 INVX1_1073 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_8173_) );
	INVX1 INVX1_1074 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_8174_) );
	NOR2X1 NOR2X1_991 ( .A(_8120_), .B(_8077_), .Y(_8175_) );
	NAND2X1 NAND2X1_1723 ( .A(_8076_), .B(_8175_), .Y(_8176_) );
	NAND2X1 NAND2X1_1724 ( .A(_8117_), .B(_8102_), .Y(_8177_) );
	OAI22X1 OAI22X1_227 ( .A(_8174_), .B(_8176_), .C(_8177_), .D(_8173_), .Y(_8178_) );
	INVX1 INVX1_1075 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_8179_) );
	INVX1 INVX1_1076 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_8180_) );
	NAND2X1 NAND2X1_1725 ( .A(_8076_), .B(_8102_), .Y(_8181_) );
	NAND2X1 NAND2X1_1726 ( .A(_8117_), .B(_8148_), .Y(_8182_) );
	OAI22X1 OAI22X1_228 ( .A(_8179_), .B(_8182_), .C(_8181_), .D(_8180_), .Y(_8183_) );
	NOR2X1 NOR2X1_992 ( .A(_8178_), .B(_8183_), .Y(_8184_) );
	INVX1 INVX1_1077 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_8185_) );
	NOR3X1 NOR3X1_700 ( .A(_8100_), .B(_8114_), .C(_8079_), .Y(_8186_) );
	NAND2X1 NAND2X1_1727 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_8186_), .Y(_8187_) );
	OR2X2 OR2X2_97 ( .A(_8112_), .B(_8094_), .Y(_8188_) );
	OAI21X1 OAI21X1_283 ( .A(_8185_), .B(_8188_), .C(_8187_), .Y(_8189_) );
	INVX1 INVX1_1078 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_8190_) );
	INVX1 INVX1_1079 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_8191_) );
	NOR2X1 NOR2X1_993 ( .A(_8120_), .B(_8090_), .Y(_8192_) );
	NAND2X1 NAND2X1_1728 ( .A(_8076_), .B(_8192_), .Y(_8193_) );
	NAND2X1 NAND2X1_1729 ( .A(_8095_), .B(_8086_), .Y(_8194_) );
	OAI22X1 OAI22X1_229 ( .A(_8193_), .B(_8191_), .C(_8190_), .D(_8194_), .Y(_8195_) );
	NOR2X1 NOR2X1_994 ( .A(_8189_), .B(_8195_), .Y(_8196_) );
	NAND3X1 NAND3X1_411 ( .A(_8172_), .B(_8196_), .C(_8184_), .Y(_8197_) );
	NOR3X1 NOR3X1_701 ( .A(_8077_), .B(_8085_), .C(_8100_), .Y(_8198_) );
	NOR3X1 NOR3X1_702 ( .A(_8094_), .B(_8120_), .C(_8084_), .Y(_8199_) );
	AOI22X1 AOI22X1_1323 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_8198_), .C(_8199_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_8200_) );
	NOR3X1 NOR3X1_703 ( .A(_8094_), .B(_8120_), .C(_8090_), .Y(_8201_) );
	NOR3X1 NOR3X1_704 ( .A(_8094_), .B(_8114_), .C(_8092_), .Y(_8202_) );
	AOI22X1 AOI22X1_1324 ( .A(_8201_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_8202_), .Y(_8203_) );
	NAND2X1 NAND2X1_1730 ( .A(_8200_), .B(_8203_), .Y(_8204_) );
	NOR3X1 NOR3X1_705 ( .A(_8092_), .B(_8077_), .C(_8104_), .Y(_8205_) );
	NOR3X1 NOR3X1_706 ( .A(_8084_), .B(_8092_), .C(_8104_), .Y(_8206_) );
	AOI22X1 AOI22X1_1325 ( .A(_8205_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_8206_), .Y(_8207_) );
	NOR3X1 NOR3X1_707 ( .A(_8075_), .B(_8120_), .C(_8084_), .Y(_8208_) );
	NOR3X1 NOR3X1_708 ( .A(_8114_), .B(_8120_), .C(_8075_), .Y(_8209_) );
	AOI22X1 AOI22X1_1326 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_8209_), .C(_8208_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_8210_) );
	NAND2X1 NAND2X1_1731 ( .A(_8210_), .B(_8207_), .Y(_8211_) );
	NOR2X1 NOR2X1_995 ( .A(_8204_), .B(_8211_), .Y(_8212_) );
	NOR3X1 NOR3X1_709 ( .A(_8100_), .B(_8120_), .C(_8084_), .Y(_8213_) );
	NOR3X1 NOR3X1_710 ( .A(_8100_), .B(_8120_), .C(_8090_), .Y(_8214_) );
	AOI22X1 AOI22X1_1327 ( .A(_8213_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_8214_), .Y(_8215_) );
	NOR3X1 NOR3X1_711 ( .A(_8100_), .B(_8114_), .C(_8092_), .Y(_8216_) );
	NOR3X1 NOR3X1_712 ( .A(_8075_), .B(_8085_), .C(_8090_), .Y(_8217_) );
	AOI22X1 AOI22X1_1328 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_8216_), .C(_8217_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_8218_) );
	NAND2X1 NAND2X1_1732 ( .A(_8215_), .B(_8218_), .Y(_8219_) );
	NOR3X1 NOR3X1_713 ( .A(_8114_), .B(_8120_), .C(_8100_), .Y(_8220_) );
	NOR3X1 NOR3X1_714 ( .A(_8090_), .B(_8085_), .C(_8104_), .Y(_8221_) );
	AOI22X1 AOI22X1_1329 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_8220_), .C(_8221_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_8222_) );
	NOR3X1 NOR3X1_715 ( .A(_8077_), .B(_8085_), .C(_8104_), .Y(_8223_) );
	NOR3X1 NOR3X1_716 ( .A(_8077_), .B(_8120_), .C(_8104_), .Y(_8224_) );
	AOI22X1 AOI22X1_1330 ( .A(_8223_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_8224_), .Y(_8225_) );
	NAND2X1 NAND2X1_1733 ( .A(_8225_), .B(_8222_), .Y(_8226_) );
	NOR2X1 NOR2X1_996 ( .A(_8219_), .B(_8226_), .Y(_8227_) );
	NAND2X1 NAND2X1_1734 ( .A(_8227_), .B(_8212_), .Y(_8228_) );
	NOR3X1 NOR3X1_717 ( .A(_8075_), .B(_8114_), .C(_8092_), .Y(_8229_) );
	NOR3X1 NOR3X1_718 ( .A(_8085_), .B(_8094_), .C(_8090_), .Y(_8230_) );
	AOI22X1 AOI22X1_1331 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_8230_), .C(_8229_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_8231_) );
	NOR3X1 NOR3X1_719 ( .A(_8079_), .B(_8077_), .C(_8104_), .Y(_8232_) );
	NOR3X1 NOR3X1_720 ( .A(_8090_), .B(_8120_), .C(_8104_), .Y(_8233_) );
	AOI22X1 AOI22X1_1332 ( .A(_8232_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_8233_), .Y(_8234_) );
	NAND2X1 NAND2X1_1735 ( .A(_8231_), .B(_8234_), .Y(_8235_) );
	NOR3X1 NOR3X1_721 ( .A(_8075_), .B(_8084_), .C(_8092_), .Y(_8236_) );
	NAND2X1 NAND2X1_1736 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_8236_), .Y(_8237_) );
	NOR3X1 NOR3X1_722 ( .A(_8094_), .B(_8114_), .C(_8079_), .Y(_8238_) );
	NAND2X1 NAND2X1_1737 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_8238_), .Y(_8239_) );
	NOR3X1 NOR3X1_723 ( .A(_8077_), .B(_8120_), .C(_8100_), .Y(_8240_) );
	NOR3X1 NOR3X1_724 ( .A(_8077_), .B(_8094_), .C(_8092_), .Y(_8241_) );
	AOI22X1 AOI22X1_1333 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_8240_), .C(_8241_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_8242_) );
	NAND3X1 NAND3X1_412 ( .A(_8237_), .B(_8239_), .C(_8242_), .Y(_8243_) );
	NOR2X1 NOR2X1_997 ( .A(_8243_), .B(_8235_), .Y(_8244_) );
	NOR3X1 NOR3X1_725 ( .A(_8077_), .B(_8100_), .C(_8092_), .Y(_8245_) );
	NOR3X1 NOR3X1_726 ( .A(_8079_), .B(_8094_), .C(_8084_), .Y(_8246_) );
	AOI22X1 AOI22X1_1334 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_8245_), .C(_8246_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_8247_) );
	NOR3X1 NOR3X1_727 ( .A(_8079_), .B(_8094_), .C(_8090_), .Y(_8248_) );
	NAND2X1 NAND2X1_1738 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_8248_), .Y(_8249_) );
	NOR3X1 NOR3X1_728 ( .A(_8084_), .B(_8085_), .C(_8104_), .Y(_8250_) );
	NAND2X1 NAND2X1_1739 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_8250_), .Y(_8251_) );
	NAND3X1 NAND3X1_413 ( .A(_8249_), .B(_8251_), .C(_8247_), .Y(_8252_) );
	NOR3X1 NOR3X1_729 ( .A(_8084_), .B(_8100_), .C(_8092_), .Y(_8253_) );
	NOR3X1 NOR3X1_730 ( .A(_8094_), .B(_8120_), .C(_8077_), .Y(_8254_) );
	AOI22X1 AOI22X1_1335 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_8254_), .C(_8253_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_8255_) );
	NOR3X1 NOR3X1_731 ( .A(_8090_), .B(_8100_), .C(_8092_), .Y(_8256_) );
	NOR3X1 NOR3X1_732 ( .A(_8094_), .B(_8114_), .C(_8085_), .Y(_8257_) );
	AOI22X1 AOI22X1_1336 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_8257_), .C(_8256_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_8258_) );
	NAND2X1 NAND2X1_1740 ( .A(_8255_), .B(_8258_), .Y(_8259_) );
	NOR2X1 NOR2X1_998 ( .A(_8259_), .B(_8252_), .Y(_8260_) );
	NAND2X1 NAND2X1_1741 ( .A(_8244_), .B(_8260_), .Y(_8261_) );
	NOR3X1 NOR3X1_733 ( .A(_8228_), .B(_8197_), .C(_8261_), .Y(_8262_) );
	INVX1 INVX1_1080 ( .A(wSelec[167]), .Y(_8263_) );
	NAND2X1 NAND2X1_1742 ( .A(wSelec[166]), .B(_8263_), .Y(_8264_) );
	INVX1 INVX1_1081 ( .A(wSelec[169]), .Y(_8265_) );
	NAND2X1 NAND2X1_1743 ( .A(wSelec[168]), .B(_8265_), .Y(_8266_) );
	NOR2X1 NOR2X1_999 ( .A(_8264_), .B(_8266_), .Y(_8267_) );
	NOR2X1 NOR2X1_1000 ( .A(wSelec[167]), .B(wSelec[166]), .Y(_8268_) );
	INVX1 INVX1_1082 ( .A(_8268_), .Y(_8269_) );
	NOR2X1 NOR2X1_1001 ( .A(_8266_), .B(_8269_), .Y(_8270_) );
	AOI22X1 AOI22X1_1337 ( .A(wData[20]), .B(_8267_), .C(_8270_), .D(wData[16]), .Y(_8271_) );
	INVX1 INVX1_1083 ( .A(wSelec[166]), .Y(_8272_) );
	NAND2X1 NAND2X1_1744 ( .A(wSelec[167]), .B(_8272_), .Y(_8273_) );
	NOR2X1 NOR2X1_1002 ( .A(_8273_), .B(_8266_), .Y(_8274_) );
	NAND2X1 NAND2X1_1745 ( .A(wData[24]), .B(_8274_), .Y(_8275_) );
	INVX1 INVX1_1084 ( .A(wSelec[168]), .Y(_8276_) );
	NAND2X1 NAND2X1_1746 ( .A(_8276_), .B(_8265_), .Y(_8277_) );
	NOR2X1 NOR2X1_1003 ( .A(_8264_), .B(_8277_), .Y(_8278_) );
	NAND2X1 NAND2X1_1747 ( .A(wSelec[167]), .B(wSelec[166]), .Y(_8279_) );
	NOR2X1 NOR2X1_1004 ( .A(_8279_), .B(_8266_), .Y(_8280_) );
	AOI22X1 AOI22X1_1338 ( .A(_8280_), .B(wData[28]), .C(wData[4]), .D(_8278_), .Y(_8281_) );
	NAND3X1 NAND3X1_414 ( .A(_8275_), .B(_8281_), .C(_8271_), .Y(_8282_) );
	NAND2X1 NAND2X1_1748 ( .A(wSelec[169]), .B(_8276_), .Y(_8283_) );
	NOR2X1 NOR2X1_1005 ( .A(_8283_), .B(_8269_), .Y(_8284_) );
	NAND2X1 NAND2X1_1749 ( .A(wData[32]), .B(_8284_), .Y(_8285_) );
	NAND2X1 NAND2X1_1750 ( .A(wSelec[168]), .B(wSelec[169]), .Y(_8286_) );
	NOR2X1 NOR2X1_1006 ( .A(_8286_), .B(_8273_), .Y(_8287_) );
	NOR2X1 NOR2X1_1007 ( .A(_8286_), .B(_8264_), .Y(_8288_) );
	AOI22X1 AOI22X1_1339 ( .A(_8287_), .B(wData[56]), .C(wData[52]), .D(_8288_), .Y(_8289_) );
	NOR2X1 NOR2X1_1008 ( .A(_8279_), .B(_8286_), .Y(_8290_) );
	NOR2X1 NOR2X1_1009 ( .A(_8279_), .B(_8283_), .Y(_8291_) );
	AOI22X1 AOI22X1_1340 ( .A(wData[60]), .B(_8290_), .C(_8291_), .D(wData[44]), .Y(_8292_) );
	NAND3X1 NAND3X1_415 ( .A(_8285_), .B(_8292_), .C(_8289_), .Y(_8293_) );
	NOR2X1 NOR2X1_1010 ( .A(_8273_), .B(_8283_), .Y(_8294_) );
	NAND2X1 NAND2X1_1751 ( .A(wData[40]), .B(_8294_), .Y(_8295_) );
	NOR2X1 NOR2X1_1011 ( .A(_8283_), .B(_8264_), .Y(_8296_) );
	NAND2X1 NAND2X1_1752 ( .A(wData[36]), .B(_8296_), .Y(_8297_) );
	NOR2X1 NOR2X1_1012 ( .A(_8277_), .B(_8269_), .Y(_8298_) );
	NAND2X1 NAND2X1_1753 ( .A(wData[0]), .B(_8298_), .Y(_8299_) );
	NAND3X1 NAND3X1_416 ( .A(_8295_), .B(_8297_), .C(_8299_), .Y(_8300_) );
	INVX1 INVX1_1085 ( .A(wData[48]), .Y(_8301_) );
	NOR2X1 NOR2X1_1013 ( .A(_8276_), .B(_8265_), .Y(_8302_) );
	NAND2X1 NAND2X1_1754 ( .A(_8268_), .B(_8302_), .Y(_8303_) );
	NOR2X1 NOR2X1_1014 ( .A(_8273_), .B(_8277_), .Y(_8304_) );
	NOR2X1 NOR2X1_1015 ( .A(_8279_), .B(_8277_), .Y(_8305_) );
	AOI22X1 AOI22X1_1341 ( .A(_8304_), .B(wData[8]), .C(wData[12]), .D(_8305_), .Y(_8306_) );
	OAI21X1 OAI21X1_284 ( .A(_8301_), .B(_8303_), .C(_8306_), .Y(_8307_) );
	OR2X2 OR2X2_98 ( .A(_8307_), .B(_8300_), .Y(_8308_) );
	NOR3X1 NOR3X1_734 ( .A(_8282_), .B(_8293_), .C(_8308_), .Y(_8309_) );
	AND2X2 AND2X2_186 ( .A(_8309_), .B(_8073_), .Y(_8310_) );
	AOI21X1 AOI21X1_201 ( .A(_8164_), .B(_8262_), .C(_8310_), .Y(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_0_) );
	INVX1 INVX1_1086 ( .A(_8181_), .Y(_8311_) );
	AOI21X1 AOI21X1_202 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_8311_), .C(_8073_), .Y(_8312_) );
	AOI22X1 AOI22X1_1342 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_8081_), .C(_8097_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_8313_) );
	AOI22X1 AOI22X1_1343 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_8101_), .C(_8107_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_8314_) );
	NAND3X1 NAND3X1_417 ( .A(_8312_), .B(_8313_), .C(_8314_), .Y(_8315_) );
	INVX1 INVX1_1087 ( .A(_8141_), .Y(_8316_) );
	AOI22X1 AOI22X1_1344 ( .A(_8166_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_8316_), .Y(_8317_) );
	AOI22X1 AOI22X1_1345 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_8240_), .C(_8119_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_8318_) );
	INVX1 INVX1_1088 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_8319_) );
	INVX1 INVX1_1089 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_8320_) );
	OAI22X1 OAI22X1_230 ( .A(_8319_), .B(_8128_), .C(_8126_), .D(_8320_), .Y(_8321_) );
	INVX1 INVX1_1090 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_8322_) );
	NAND2X1 NAND2X1_1755 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_8229_), .Y(_8323_) );
	OAI21X1 OAI21X1_285 ( .A(_8322_), .B(_8134_), .C(_8323_), .Y(_8324_) );
	NOR2X1 NOR2X1_1016 ( .A(_8321_), .B(_8324_), .Y(_8325_) );
	NAND3X1 NAND3X1_418 ( .A(_8317_), .B(_8318_), .C(_8325_), .Y(_8326_) );
	INVX1 INVX1_1091 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_8327_) );
	NAND2X1 NAND2X1_1756 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_8113_), .Y(_8328_) );
	OAI21X1 OAI21X1_286 ( .A(_8327_), .B(_8143_), .C(_8328_), .Y(_8329_) );
	INVX1 INVX1_1092 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_8330_) );
	INVX1 INVX1_1093 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_8331_) );
	OAI22X1 OAI22X1_231 ( .A(_8330_), .B(_8149_), .C(_8147_), .D(_8331_), .Y(_8332_) );
	NOR2X1 NOR2X1_1017 ( .A(_8332_), .B(_8329_), .Y(_8333_) );
	AOI22X1 AOI22X1_1346 ( .A(_8233_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_8206_), .Y(_8334_) );
	AND2X2 AND2X2_187 ( .A(_8080_), .B(_8095_), .Y(_8335_) );
	AOI22X1 AOI22X1_1347 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_8205_), .C(_8335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_8336_) );
	NAND3X1 NAND3X1_419 ( .A(_8334_), .B(_8336_), .C(_8333_), .Y(_8337_) );
	NOR3X1 NOR3X1_735 ( .A(_8337_), .B(_8315_), .C(_8326_), .Y(_8338_) );
	INVX1 INVX1_1094 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_8339_) );
	NAND2X1 NAND2X1_1757 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_8168_), .Y(_8340_) );
	OAI21X1 OAI21X1_287 ( .A(_8170_), .B(_8339_), .C(_8340_), .Y(_8341_) );
	AOI21X1 AOI21X1_203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_8217_), .C(_8341_), .Y(_8342_) );
	INVX1 INVX1_1095 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_8343_) );
	INVX1 INVX1_1096 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_8344_) );
	OAI22X1 OAI22X1_232 ( .A(_8344_), .B(_8176_), .C(_8177_), .D(_8343_), .Y(_8345_) );
	INVX1 INVX1_1097 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_8346_) );
	NAND2X1 NAND2X1_1758 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_8186_), .Y(_8347_) );
	OAI21X1 OAI21X1_288 ( .A(_8087_), .B(_8346_), .C(_8347_), .Y(_8348_) );
	NOR2X1 NOR2X1_1018 ( .A(_8348_), .B(_8345_), .Y(_8349_) );
	INVX1 INVX1_1098 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_8350_) );
	INVX1 INVX1_1099 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_8351_) );
	OAI22X1 OAI22X1_233 ( .A(_8182_), .B(_8351_), .C(_8188_), .D(_8350_), .Y(_8352_) );
	INVX1 INVX1_1100 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_8353_) );
	NOR2X1 NOR2X1_1019 ( .A(_8353_), .B(_8193_), .Y(_8354_) );
	INVX1 INVX1_1101 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_8355_) );
	NOR2X1 NOR2X1_1020 ( .A(_8355_), .B(_8194_), .Y(_8356_) );
	NOR3X1 NOR3X1_736 ( .A(_8354_), .B(_8352_), .C(_8356_), .Y(_8357_) );
	NAND3X1 NAND3X1_420 ( .A(_8349_), .B(_8342_), .C(_8357_), .Y(_8358_) );
	AOI22X1 AOI22X1_1348 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_8198_), .C(_8199_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_8359_) );
	AOI22X1 AOI22X1_1349 ( .A(_8201_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_8202_), .Y(_8360_) );
	NAND2X1 NAND2X1_1759 ( .A(_8359_), .B(_8360_), .Y(_8361_) );
	AOI22X1 AOI22X1_1350 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_8209_), .C(_8208_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_8362_) );
	AOI22X1 AOI22X1_1351 ( .A(_8152_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_8159_), .Y(_8363_) );
	NAND2X1 NAND2X1_1760 ( .A(_8362_), .B(_8363_), .Y(_8364_) );
	NOR2X1 NOR2X1_1021 ( .A(_8361_), .B(_8364_), .Y(_8365_) );
	AOI22X1 AOI22X1_1352 ( .A(_8213_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_8214_), .Y(_8366_) );
	AOI22X1 AOI22X1_1353 ( .A(_8115_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_8216_), .Y(_8367_) );
	NAND2X1 NAND2X1_1761 ( .A(_8366_), .B(_8367_), .Y(_8368_) );
	AOI22X1 AOI22X1_1354 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_8220_), .C(_8221_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_8369_) );
	AOI22X1 AOI22X1_1355 ( .A(_8223_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_8224_), .Y(_8370_) );
	NAND2X1 NAND2X1_1762 ( .A(_8370_), .B(_8369_), .Y(_8371_) );
	NOR2X1 NOR2X1_1022 ( .A(_8368_), .B(_8371_), .Y(_8372_) );
	NAND2X1 NAND2X1_1763 ( .A(_8372_), .B(_8365_), .Y(_8373_) );
	AOI22X1 AOI22X1_1356 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_8230_), .C(_8131_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_8374_) );
	AOI22X1 AOI22X1_1357 ( .A(_8154_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_8232_), .Y(_8375_) );
	NAND2X1 NAND2X1_1764 ( .A(_8374_), .B(_8375_), .Y(_8376_) );
	AOI22X1 AOI22X1_1358 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_8121_), .C(_8241_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_8377_) );
	NAND2X1 NAND2X1_1765 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_8236_), .Y(_8378_) );
	NAND2X1 NAND2X1_1766 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_8238_), .Y(_8379_) );
	NAND3X1 NAND3X1_421 ( .A(_8378_), .B(_8379_), .C(_8377_), .Y(_8380_) );
	NOR2X1 NOR2X1_1023 ( .A(_8380_), .B(_8376_), .Y(_8381_) );
	AOI22X1 AOI22X1_1359 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_8245_), .C(_8246_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_8382_) );
	NAND2X1 NAND2X1_1767 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_8248_), .Y(_8383_) );
	NAND2X1 NAND2X1_1768 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_8250_), .Y(_8384_) );
	NAND3X1 NAND3X1_422 ( .A(_8383_), .B(_8384_), .C(_8382_), .Y(_8385_) );
	AOI22X1 AOI22X1_1360 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_8254_), .C(_8253_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_8386_) );
	AOI22X1 AOI22X1_1361 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_8257_), .C(_8256_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_8387_) );
	NAND2X1 NAND2X1_1769 ( .A(_8386_), .B(_8387_), .Y(_8388_) );
	NOR2X1 NOR2X1_1024 ( .A(_8388_), .B(_8385_), .Y(_8389_) );
	NAND2X1 NAND2X1_1770 ( .A(_8381_), .B(_8389_), .Y(_8390_) );
	NOR3X1 NOR3X1_737 ( .A(_8373_), .B(_8358_), .C(_8390_), .Y(_8391_) );
	AOI21X1 AOI21X1_204 ( .A(wData[21]), .B(_8267_), .C(_8072_), .Y(_8392_) );
	AOI22X1 AOI22X1_1362 ( .A(_8270_), .B(wData[17]), .C(wData[1]), .D(_8298_), .Y(_8393_) );
	AOI22X1 AOI22X1_1363 ( .A(_8291_), .B(wData[45]), .C(wData[25]), .D(_8274_), .Y(_8394_) );
	NAND3X1 NAND3X1_423 ( .A(_8392_), .B(_8394_), .C(_8393_), .Y(_8395_) );
	NAND3X1 NAND3X1_424 ( .A(wData[49]), .B(_8268_), .C(_8302_), .Y(_8396_) );
	AOI22X1 AOI22X1_1364 ( .A(wData[61]), .B(_8290_), .C(_8278_), .D(wData[5]), .Y(_8397_) );
	AND2X2 AND2X2_188 ( .A(_8397_), .B(_8396_), .Y(_8398_) );
	AOI22X1 AOI22X1_1365 ( .A(_8287_), .B(wData[57]), .C(wData[41]), .D(_8294_), .Y(_8399_) );
	AOI22X1 AOI22X1_1366 ( .A(wData[53]), .B(_8288_), .C(_8284_), .D(wData[33]), .Y(_8400_) );
	AND2X2 AND2X2_189 ( .A(_8400_), .B(_8399_), .Y(_8401_) );
	AOI22X1 AOI22X1_1367 ( .A(_8304_), .B(wData[9]), .C(wData[13]), .D(_8305_), .Y(_8402_) );
	AOI22X1 AOI22X1_1368 ( .A(_8280_), .B(wData[29]), .C(wData[37]), .D(_8296_), .Y(_8403_) );
	AND2X2 AND2X2_190 ( .A(_8402_), .B(_8403_), .Y(_8404_) );
	NAND3X1 NAND3X1_425 ( .A(_8398_), .B(_8404_), .C(_8401_), .Y(_8405_) );
	NOR2X1 NOR2X1_1025 ( .A(_8395_), .B(_8405_), .Y(_8406_) );
	AOI21X1 AOI21X1_205 ( .A(_8338_), .B(_8391_), .C(_8406_), .Y(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_1_) );
	AOI21X1 AOI21X1_206 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_8311_), .C(_8073_), .Y(_8407_) );
	INVX1 INVX1_1102 ( .A(_8170_), .Y(_8408_) );
	AOI22X1 AOI22X1_1369 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_8081_), .C(_8408_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_8409_) );
	INVX1 INVX1_1103 ( .A(_8182_), .Y(_8410_) );
	AOI22X1 AOI22X1_1370 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_8217_), .C(_8410_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_8411_) );
	NAND3X1 NAND3X1_426 ( .A(_8411_), .B(_8407_), .C(_8409_), .Y(_8412_) );
	AOI22X1 AOI22X1_1371 ( .A(_8166_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_8316_), .Y(_8413_) );
	AOI22X1 AOI22X1_1372 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_8115_), .C(_8088_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_8414_) );
	INVX1 INVX1_1104 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_8415_) );
	NAND2X1 NAND2X1_1771 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_8205_), .Y(_8416_) );
	OAI21X1 OAI21X1_289 ( .A(_8415_), .B(_8177_), .C(_8416_), .Y(_8417_) );
	INVX1 INVX1_1105 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_8418_) );
	NAND2X1 NAND2X1_1772 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_8131_), .Y(_8419_) );
	OAI21X1 OAI21X1_290 ( .A(_8418_), .B(_8134_), .C(_8419_), .Y(_8420_) );
	NOR2X1 NOR2X1_1026 ( .A(_8417_), .B(_8420_), .Y(_8421_) );
	NAND3X1 NAND3X1_427 ( .A(_8413_), .B(_8414_), .C(_8421_), .Y(_8422_) );
	INVX1 INVX1_1106 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_8423_) );
	NAND2X1 NAND2X1_1773 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_8113_), .Y(_8424_) );
	OAI21X1 OAI21X1_291 ( .A(_8423_), .B(_8143_), .C(_8424_), .Y(_8425_) );
	INVX1 INVX1_1107 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_8426_) );
	INVX1 INVX1_1108 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_8427_) );
	OAI22X1 OAI22X1_234 ( .A(_8426_), .B(_8149_), .C(_8147_), .D(_8427_), .Y(_8428_) );
	NOR2X1 NOR2X1_1027 ( .A(_8428_), .B(_8425_), .Y(_8429_) );
	AOI22X1 AOI22X1_1373 ( .A(_8233_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_8206_), .Y(_8430_) );
	AND2X2 AND2X2_191 ( .A(_8105_), .B(_8127_), .Y(_8431_) );
	AOI22X1 AOI22X1_1374 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_8431_), .C(_8335_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_8432_) );
	NAND3X1 NAND3X1_428 ( .A(_8430_), .B(_8432_), .C(_8429_), .Y(_8433_) );
	NOR3X1 NOR3X1_738 ( .A(_8433_), .B(_8412_), .C(_8422_), .Y(_8434_) );
	INVX1 INVX1_1109 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_8435_) );
	NOR3X1 NOR3X1_739 ( .A(_8435_), .B(_8100_), .C(_8099_), .Y(_8436_) );
	AND2X2 AND2X2_192 ( .A(_8121_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_8437_) );
	AND2X2 AND2X2_193 ( .A(_8241_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_8438_) );
	NOR3X1 NOR3X1_740 ( .A(_8438_), .B(_8437_), .C(_8436_), .Y(_8439_) );
	INVX1 INVX1_1110 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_8440_) );
	INVX1 INVX1_1111 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_8441_) );
	OAI22X1 OAI22X1_235 ( .A(_8441_), .B(_8176_), .C(_8126_), .D(_8440_), .Y(_8442_) );
	INVX1 INVX1_1112 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_8443_) );
	INVX1 INVX1_1113 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_8444_) );
	NAND2X1 NAND2X1_1774 ( .A(_8117_), .B(_8118_), .Y(_8445_) );
	OAI22X1 OAI22X1_236 ( .A(_8445_), .B(_8444_), .C(_8443_), .D(_8096_), .Y(_8446_) );
	NOR2X1 NOR2X1_1028 ( .A(_8442_), .B(_8446_), .Y(_8447_) );
	INVX1 INVX1_1114 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_8448_) );
	NOR3X1 NOR3X1_741 ( .A(_8077_), .B(_8094_), .C(_8085_), .Y(_8449_) );
	NAND2X1 NAND2X1_1775 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_8449_), .Y(_8450_) );
	OAI21X1 OAI21X1_292 ( .A(_8106_), .B(_8448_), .C(_8450_), .Y(_8451_) );
	INVX1 INVX1_1115 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_8452_) );
	INVX1 INVX1_1116 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_8453_) );
	OAI22X1 OAI22X1_237 ( .A(_8193_), .B(_8453_), .C(_8452_), .D(_8194_), .Y(_8454_) );
	NOR2X1 NOR2X1_1029 ( .A(_8451_), .B(_8454_), .Y(_8455_) );
	NAND3X1 NAND3X1_429 ( .A(_8439_), .B(_8455_), .C(_8447_), .Y(_8456_) );
	AOI22X1 AOI22X1_1375 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_8198_), .C(_8199_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_8457_) );
	AOI22X1 AOI22X1_1376 ( .A(_8201_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_8202_), .Y(_8458_) );
	NAND2X1 NAND2X1_1776 ( .A(_8457_), .B(_8458_), .Y(_8459_) );
	AOI22X1 AOI22X1_1377 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_8209_), .C(_8208_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_8460_) );
	AOI22X1 AOI22X1_1378 ( .A(_8152_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_8159_), .Y(_8461_) );
	NAND2X1 NAND2X1_1777 ( .A(_8460_), .B(_8461_), .Y(_8462_) );
	NOR2X1 NOR2X1_1030 ( .A(_8459_), .B(_8462_), .Y(_8463_) );
	AOI22X1 AOI22X1_1379 ( .A(_8213_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_8214_), .Y(_8464_) );
	AOI22X1 AOI22X1_1380 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_8240_), .C(_8216_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_8465_) );
	NAND2X1 NAND2X1_1778 ( .A(_8465_), .B(_8464_), .Y(_8466_) );
	AOI22X1 AOI22X1_1381 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_8220_), .C(_8221_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_8467_) );
	AOI22X1 AOI22X1_1382 ( .A(_8223_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_8224_), .Y(_8468_) );
	NAND2X1 NAND2X1_1779 ( .A(_8468_), .B(_8467_), .Y(_8469_) );
	NOR2X1 NOR2X1_1031 ( .A(_8466_), .B(_8469_), .Y(_8470_) );
	NAND2X1 NAND2X1_1780 ( .A(_8470_), .B(_8463_), .Y(_8471_) );
	AOI22X1 AOI22X1_1383 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_8230_), .C(_8229_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_8472_) );
	AOI22X1 AOI22X1_1384 ( .A(_8154_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_8232_), .Y(_8473_) );
	NAND2X1 NAND2X1_1781 ( .A(_8472_), .B(_8473_), .Y(_8474_) );
	AOI22X1 AOI22X1_1385 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_8238_), .C(_8236_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_8475_) );
	AOI22X1 AOI22X1_1386 ( .A(_8168_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_8186_), .Y(_8476_) );
	NAND2X1 NAND2X1_1782 ( .A(_8476_), .B(_8475_), .Y(_8477_) );
	NOR2X1 NOR2X1_1032 ( .A(_8477_), .B(_8474_), .Y(_8478_) );
	AOI22X1 AOI22X1_1387 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_8245_), .C(_8246_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_8479_) );
	NAND2X1 NAND2X1_1783 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_8248_), .Y(_8480_) );
	NAND2X1 NAND2X1_1784 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_8250_), .Y(_8481_) );
	NAND3X1 NAND3X1_430 ( .A(_8480_), .B(_8481_), .C(_8479_), .Y(_8482_) );
	AOI22X1 AOI22X1_1388 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_8254_), .C(_8253_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_8483_) );
	AOI22X1 AOI22X1_1389 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_8257_), .C(_8256_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_8484_) );
	NAND2X1 NAND2X1_1785 ( .A(_8483_), .B(_8484_), .Y(_8485_) );
	NOR2X1 NOR2X1_1033 ( .A(_8485_), .B(_8482_), .Y(_8486_) );
	NAND2X1 NAND2X1_1786 ( .A(_8478_), .B(_8486_), .Y(_8487_) );
	NOR3X1 NOR3X1_742 ( .A(_8471_), .B(_8456_), .C(_8487_), .Y(_8488_) );
	AOI22X1 AOI22X1_1390 ( .A(_8294_), .B(wData[42]), .C(wData[38]), .D(_8296_), .Y(_8489_) );
	AOI22X1 AOI22X1_1391 ( .A(_8291_), .B(wData[46]), .C(_8298_), .D(wData[2]), .Y(_8490_) );
	NAND2X1 NAND2X1_1787 ( .A(_8489_), .B(_8490_), .Y(_8491_) );
	AOI21X1 AOI21X1_207 ( .A(wData[34]), .B(_8284_), .C(_8491_), .Y(_8492_) );
	INVX1 INVX1_1117 ( .A(wData[50]), .Y(_8493_) );
	AOI22X1 AOI22X1_1392 ( .A(_8304_), .B(wData[10]), .C(wData[14]), .D(_8305_), .Y(_8494_) );
	OAI21X1 OAI21X1_293 ( .A(_8493_), .B(_8303_), .C(_8494_), .Y(_8495_) );
	AOI22X1 AOI22X1_1393 ( .A(_8267_), .B(wData[22]), .C(wData[18]), .D(_8270_), .Y(_8496_) );
	NAND2X1 NAND2X1_1788 ( .A(wData[26]), .B(_8274_), .Y(_8497_) );
	AOI22X1 AOI22X1_1394 ( .A(_8280_), .B(wData[30]), .C(wData[6]), .D(_8278_), .Y(_8498_) );
	NAND3X1 NAND3X1_431 ( .A(_8497_), .B(_8498_), .C(_8496_), .Y(_8499_) );
	NOR2X1 NOR2X1_1034 ( .A(_8495_), .B(_8499_), .Y(_8500_) );
	NAND2X1 NAND2X1_1789 ( .A(wData[58]), .B(_8287_), .Y(_8501_) );
	NAND2X1 NAND2X1_1790 ( .A(wData[54]), .B(_8288_), .Y(_8502_) );
	NAND2X1 NAND2X1_1791 ( .A(_8501_), .B(_8502_), .Y(_8503_) );
	AOI21X1 AOI21X1_208 ( .A(wData[62]), .B(_8290_), .C(_8503_), .Y(_8504_) );
	NAND3X1 NAND3X1_432 ( .A(_8492_), .B(_8504_), .C(_8500_), .Y(_8505_) );
	NOR2X1 NOR2X1_1035 ( .A(_8072_), .B(_8505_), .Y(_8506_) );
	AOI21X1 AOI21X1_209 ( .A(_8434_), .B(_8488_), .C(_8506_), .Y(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_2_) );
	AOI21X1 AOI21X1_210 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_8316_), .C(_8073_), .Y(_8507_) );
	AOI22X1 AOI22X1_1395 ( .A(_8088_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_8408_), .Y(_8508_) );
	AOI22X1 AOI22X1_1396 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_8410_), .C(_8166_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_8509_) );
	NAND3X1 NAND3X1_433 ( .A(_8509_), .B(_8507_), .C(_8508_), .Y(_8510_) );
	AOI22X1 AOI22X1_1397 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_8115_), .C(_8113_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_8511_) );
	AOI22X1 AOI22X1_1398 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_8186_), .C(_8311_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_8512_) );
	INVX1 INVX1_1118 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_8513_) );
	INVX1 INVX1_1119 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_8514_) );
	OAI22X1 OAI22X1_238 ( .A(_8513_), .B(_8128_), .C(_8177_), .D(_8514_), .Y(_8515_) );
	INVX1 INVX1_1120 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_8516_) );
	NAND2X1 NAND2X1_1792 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_8229_), .Y(_8517_) );
	OAI21X1 OAI21X1_294 ( .A(_8516_), .B(_8134_), .C(_8517_), .Y(_8518_) );
	NOR2X1 NOR2X1_1036 ( .A(_8515_), .B(_8518_), .Y(_8519_) );
	NAND3X1 NAND3X1_434 ( .A(_8511_), .B(_8512_), .C(_8519_), .Y(_8520_) );
	AND2X2 AND2X2_194 ( .A(_8142_), .B(_8076_), .Y(_8521_) );
	AOI22X1 AOI22X1_1399 ( .A(_8081_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_8521_), .Y(_8522_) );
	AND2X2 AND2X2_195 ( .A(_8140_), .B(_8105_), .Y(_8523_) );
	AND2X2 AND2X2_196 ( .A(_8148_), .B(_8105_), .Y(_8524_) );
	AOI22X1 AOI22X1_1400 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_8524_), .C(_8523_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_8525_) );
	NAND2X1 NAND2X1_1793 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_8233_), .Y(_8526_) );
	NAND2X1 NAND2X1_1794 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_8206_), .Y(_8527_) );
	NAND2X1 NAND2X1_1795 ( .A(_8526_), .B(_8527_), .Y(_8528_) );
	INVX1 INVX1_1121 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_8529_) );
	NAND2X1 NAND2X1_1796 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_8205_), .Y(_8530_) );
	OAI21X1 OAI21X1_295 ( .A(_8529_), .B(_8158_), .C(_8530_), .Y(_8531_) );
	NOR2X1 NOR2X1_1037 ( .A(_8528_), .B(_8531_), .Y(_8532_) );
	NAND3X1 NAND3X1_435 ( .A(_8522_), .B(_8525_), .C(_8532_), .Y(_8533_) );
	NOR3X1 NOR3X1_743 ( .A(_8520_), .B(_8510_), .C(_8533_), .Y(_8534_) );
	INVX1 INVX1_1122 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_8535_) );
	NAND2X1 NAND2X1_1797 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_8121_), .Y(_8536_) );
	OAI21X1 OAI21X1_296 ( .A(_8126_), .B(_8535_), .C(_8536_), .Y(_8537_) );
	AOI21X1 AOI21X1_211 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_8101_), .C(_8537_), .Y(_8538_) );
	INVX1 INVX1_1123 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_8539_) );
	INVX1 INVX1_1124 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_8540_) );
	OAI22X1 OAI22X1_239 ( .A(_8445_), .B(_8540_), .C(_8539_), .D(_8096_), .Y(_8541_) );
	INVX1 INVX1_1125 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_8542_) );
	NAND2X1 NAND2X1_1798 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_8241_), .Y(_8543_) );
	OAI21X1 OAI21X1_297 ( .A(_8106_), .B(_8542_), .C(_8543_), .Y(_8544_) );
	NOR2X1 NOR2X1_1038 ( .A(_8544_), .B(_8541_), .Y(_8545_) );
	INVX1 INVX1_1126 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_8546_) );
	INVX1 INVX1_1127 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_8547_) );
	OAI22X1 OAI22X1_240 ( .A(_8193_), .B(_8547_), .C(_8546_), .D(_8194_), .Y(_8548_) );
	INVX1 INVX1_1128 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_8549_) );
	NAND2X1 NAND2X1_1799 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_8240_), .Y(_8550_) );
	OAI21X1 OAI21X1_298 ( .A(_8549_), .B(_8176_), .C(_8550_), .Y(_8551_) );
	NOR2X1 NOR2X1_1039 ( .A(_8551_), .B(_8548_), .Y(_8552_) );
	NAND3X1 NAND3X1_436 ( .A(_8538_), .B(_8552_), .C(_8545_), .Y(_8553_) );
	AOI22X1 AOI22X1_1401 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_8198_), .C(_8199_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_8554_) );
	AOI22X1 AOI22X1_1402 ( .A(_8201_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_8202_), .Y(_8555_) );
	NAND2X1 NAND2X1_1800 ( .A(_8554_), .B(_8555_), .Y(_8556_) );
	AOI22X1 AOI22X1_1403 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_8209_), .C(_8208_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_8557_) );
	AOI22X1 AOI22X1_1404 ( .A(_8152_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_8159_), .Y(_8558_) );
	NAND2X1 NAND2X1_1801 ( .A(_8557_), .B(_8558_), .Y(_8559_) );
	NOR2X1 NOR2X1_1040 ( .A(_8556_), .B(_8559_), .Y(_8560_) );
	AOI22X1 AOI22X1_1405 ( .A(_8213_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_8214_), .Y(_8561_) );
	AOI22X1 AOI22X1_1406 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_8449_), .C(_8216_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_8562_) );
	NAND2X1 NAND2X1_1802 ( .A(_8562_), .B(_8561_), .Y(_8563_) );
	AOI22X1 AOI22X1_1407 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_8220_), .C(_8221_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_8564_) );
	AOI22X1 AOI22X1_1408 ( .A(_8223_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_8224_), .Y(_8565_) );
	NAND2X1 NAND2X1_1803 ( .A(_8565_), .B(_8564_), .Y(_8566_) );
	NOR2X1 NOR2X1_1041 ( .A(_8563_), .B(_8566_), .Y(_8567_) );
	NAND2X1 NAND2X1_1804 ( .A(_8567_), .B(_8560_), .Y(_8568_) );
	AOI22X1 AOI22X1_1409 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_8230_), .C(_8131_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_8569_) );
	AOI22X1 AOI22X1_1410 ( .A(_8154_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_8232_), .Y(_8570_) );
	NAND2X1 NAND2X1_1805 ( .A(_8569_), .B(_8570_), .Y(_8571_) );
	AOI22X1 AOI22X1_1411 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_8238_), .C(_8236_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_8572_) );
	AOI22X1 AOI22X1_1412 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_8168_), .C(_8217_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_8573_) );
	NAND2X1 NAND2X1_1806 ( .A(_8573_), .B(_8572_), .Y(_8574_) );
	NOR2X1 NOR2X1_1042 ( .A(_8574_), .B(_8571_), .Y(_8575_) );
	AOI22X1 AOI22X1_1413 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_8245_), .C(_8246_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_8576_) );
	NAND2X1 NAND2X1_1807 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_8248_), .Y(_8577_) );
	NAND2X1 NAND2X1_1808 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_8250_), .Y(_8578_) );
	NAND3X1 NAND3X1_437 ( .A(_8577_), .B(_8578_), .C(_8576_), .Y(_8579_) );
	AOI22X1 AOI22X1_1414 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_8254_), .C(_8253_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_8580_) );
	AOI22X1 AOI22X1_1415 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_8257_), .C(_8256_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_8581_) );
	NAND2X1 NAND2X1_1809 ( .A(_8580_), .B(_8581_), .Y(_8582_) );
	NOR2X1 NOR2X1_1043 ( .A(_8582_), .B(_8579_), .Y(_8583_) );
	NAND2X1 NAND2X1_1810 ( .A(_8575_), .B(_8583_), .Y(_8584_) );
	NOR3X1 NOR3X1_744 ( .A(_8568_), .B(_8553_), .C(_8584_), .Y(_8585_) );
	NAND2X1 NAND2X1_1811 ( .A(wData[59]), .B(_8287_), .Y(_8586_) );
	OAI21X1 OAI21X1_299 ( .A(_8071_), .B(wBusy_bF_buf1), .C(_8586_), .Y(_8587_) );
	NAND2X1 NAND2X1_1812 ( .A(wData[7]), .B(_8278_), .Y(_8588_) );
	NAND2X1 NAND2X1_1813 ( .A(wData[55]), .B(_8288_), .Y(_8589_) );
	AOI22X1 AOI22X1_1416 ( .A(wData[63]), .B(_8290_), .C(_8280_), .D(wData[31]), .Y(_8590_) );
	NAND3X1 NAND3X1_438 ( .A(_8588_), .B(_8589_), .C(_8590_), .Y(_8591_) );
	OR2X2 OR2X2_99 ( .A(_8591_), .B(_8587_), .Y(_8592_) );
	INVX1 INVX1_1129 ( .A(wData[51]), .Y(_8593_) );
	NAND2X1 NAND2X1_1814 ( .A(wData[47]), .B(_8291_), .Y(_8594_) );
	OAI21X1 OAI21X1_300 ( .A(_8593_), .B(_8303_), .C(_8594_), .Y(_8595_) );
	AOI21X1 AOI21X1_212 ( .A(wData[3]), .B(_8298_), .C(_8595_), .Y(_8596_) );
	AOI22X1 AOI22X1_1417 ( .A(_8304_), .B(wData[11]), .C(wData[15]), .D(_8305_), .Y(_8597_) );
	AOI22X1 AOI22X1_1418 ( .A(_8267_), .B(wData[23]), .C(wData[27]), .D(_8274_), .Y(_8598_) );
	AND2X2 AND2X2_197 ( .A(_8597_), .B(_8598_), .Y(_8599_) );
	NAND2X1 NAND2X1_1815 ( .A(wData[39]), .B(_8296_), .Y(_8600_) );
	NAND2X1 NAND2X1_1816 ( .A(wData[43]), .B(_8294_), .Y(_8601_) );
	NAND2X1 NAND2X1_1817 ( .A(_8600_), .B(_8601_), .Y(_8602_) );
	NAND2X1 NAND2X1_1818 ( .A(wData[19]), .B(_8270_), .Y(_8603_) );
	NAND2X1 NAND2X1_1819 ( .A(wData[35]), .B(_8284_), .Y(_8604_) );
	NAND2X1 NAND2X1_1820 ( .A(_8603_), .B(_8604_), .Y(_8605_) );
	NOR2X1 NOR2X1_1044 ( .A(_8602_), .B(_8605_), .Y(_8606_) );
	NAND3X1 NAND3X1_439 ( .A(_8599_), .B(_8596_), .C(_8606_), .Y(_8607_) );
	NOR2X1 NOR2X1_1045 ( .A(_8592_), .B(_8607_), .Y(_8608_) );
	AOI21X1 AOI21X1_213 ( .A(_8534_), .B(_8585_), .C(_8608_), .Y(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_3_) );
	NOR2X1 NOR2X1_1046 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(scheduler_block_scheduler_ctr_1_bF_buf5), .Y(_8699_) );
	OAI21X1 OAI21X1_301 ( .A(_8699_), .B(rst_bF_buf3), .C(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_0_), .Y(_8700_) );
	INVX4 INVX4_1 ( .A(rst_bF_buf2), .Y(_8701_) );
	INVX4 INVX4_2 ( .A(scheduler_block_scheduler_ctr_1_bF_buf4), .Y(_8702_) );
	NAND3X1 NAND3X1_440 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_0_), .C(_8702_), .Y(_8703_) );
	NAND3X1 NAND3X1_441 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(scheduler_block_scheduler_ctr_1_bF_buf3), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_0_), .Y(_8704_) );
	INVX4 INVX4_3 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .Y(_8705_) );
	NAND3X1 NAND3X1_442 ( .A(scheduler_block_scheduler_ctr_1_bF_buf2), .B(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_0_), .C(_8705_), .Y(_8706_) );
	NAND3X1 NAND3X1_443 ( .A(_8704_), .B(_8703_), .C(_8706_), .Y(_8707_) );
	NAND2X1 NAND2X1_1821 ( .A(_8701__bF_buf3), .B(_8707_), .Y(_8708_) );
	NAND2X1 NAND2X1_1822 ( .A(_8700_), .B(_8708_), .Y(_8610__0_) );
	OAI21X1 OAI21X1_302 ( .A(_8699_), .B(rst_bF_buf1), .C(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_1_), .Y(_8709_) );
	NAND3X1 NAND3X1_444 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_1_), .C(_8702_), .Y(_8710_) );
	NAND3X1 NAND3X1_445 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf1), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_1_), .Y(_8711_) );
	NAND3X1 NAND3X1_446 ( .A(scheduler_block_scheduler_ctr_1_bF_buf0), .B(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_1_), .C(_8705_), .Y(_8611_) );
	NAND3X1 NAND3X1_447 ( .A(_8711_), .B(_8710_), .C(_8611_), .Y(_8612_) );
	NAND2X1 NAND2X1_1823 ( .A(_8701__bF_buf2), .B(_8612_), .Y(_8613_) );
	NAND2X1 NAND2X1_1824 ( .A(_8709_), .B(_8613_), .Y(_8610__1_) );
	OAI21X1 OAI21X1_303 ( .A(_8699_), .B(rst_bF_buf0), .C(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_2_), .Y(_8614_) );
	NAND3X1 NAND3X1_448 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_2_), .C(_8702_), .Y(_8615_) );
	NAND3X1 NAND3X1_449 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(scheduler_block_scheduler_ctr_1_bF_buf5), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_2_), .Y(_8616_) );
	NAND3X1 NAND3X1_450 ( .A(scheduler_block_scheduler_ctr_1_bF_buf4), .B(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_2_), .C(_8705_), .Y(_8617_) );
	NAND3X1 NAND3X1_451 ( .A(_8616_), .B(_8615_), .C(_8617_), .Y(_8618_) );
	NAND2X1 NAND2X1_1825 ( .A(_8701__bF_buf1), .B(_8618_), .Y(_8619_) );
	NAND2X1 NAND2X1_1826 ( .A(_8614_), .B(_8619_), .Y(_8610__2_) );
	OAI21X1 OAI21X1_304 ( .A(_8699_), .B(rst_bF_buf3), .C(input_selector_block_input_selector_i_3__input_selector_j_0__input_selector_r_3_), .Y(_8620_) );
	NAND3X1 NAND3X1_452 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(input_selector_block_input_selector_i_2__input_selector_j_0__input_selector_r_3_), .C(_8702_), .Y(_8621_) );
	NAND3X1 NAND3X1_453 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .B(scheduler_block_scheduler_ctr_1_bF_buf3), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_3_), .Y(_8622_) );
	NAND3X1 NAND3X1_454 ( .A(scheduler_block_scheduler_ctr_1_bF_buf2), .B(input_selector_block_input_selector_i_1__input_selector_j_0__input_selector_r_3_), .C(_8705_), .Y(_8623_) );
	NAND3X1 NAND3X1_455 ( .A(_8622_), .B(_8621_), .C(_8623_), .Y(_8624_) );
	NAND2X1 NAND2X1_1827 ( .A(_8701__bF_buf0), .B(_8624_), .Y(_8625_) );
	NAND2X1 NAND2X1_1828 ( .A(_8620_), .B(_8625_), .Y(_8610__3_) );
	OAI21X1 OAI21X1_305 ( .A(_8699_), .B(rst_bF_buf2), .C(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_0_), .Y(_8626_) );
	NAND3X1 NAND3X1_456 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_0_), .C(_8702_), .Y(_8627_) );
	NAND3X1 NAND3X1_457 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf1), .C(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_0_), .Y(_8628_) );
	NAND3X1 NAND3X1_458 ( .A(scheduler_block_scheduler_ctr_1_bF_buf0), .B(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_0_), .C(_8705_), .Y(_8629_) );
	NAND3X1 NAND3X1_459 ( .A(_8628_), .B(_8627_), .C(_8629_), .Y(_8630_) );
	NAND2X1 NAND2X1_1829 ( .A(_8701__bF_buf3), .B(_8630_), .Y(_8631_) );
	NAND2X1 NAND2X1_1830 ( .A(_8626_), .B(_8631_), .Y(_8610__4_) );
	OAI21X1 OAI21X1_306 ( .A(_8699_), .B(rst_bF_buf1), .C(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_1_), .Y(_8632_) );
	NAND3X1 NAND3X1_460 ( .A(scheduler_block_scheduler_ctr_1_bF_buf5), .B(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_1_), .C(_8705_), .Y(_8633_) );
	NAND3X1 NAND3X1_461 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_1_), .C(_8702_), .Y(_8634_) );
	NAND3X1 NAND3X1_462 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(scheduler_block_scheduler_ctr_1_bF_buf4), .C(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_1_), .Y(_8635_) );
	NAND3X1 NAND3X1_463 ( .A(_8635_), .B(_8633_), .C(_8634_), .Y(_8636_) );
	NAND2X1 NAND2X1_1831 ( .A(_8701__bF_buf2), .B(_8636_), .Y(_8637_) );
	NAND2X1 NAND2X1_1832 ( .A(_8632_), .B(_8637_), .Y(_8610__5_) );
	OAI21X1 OAI21X1_307 ( .A(_8699_), .B(rst_bF_buf0), .C(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_2_), .Y(_8638_) );
	NAND3X1 NAND3X1_464 ( .A(scheduler_block_scheduler_ctr_1_bF_buf3), .B(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_2_), .C(_8705_), .Y(_8639_) );
	NAND3X1 NAND3X1_465 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_2_), .C(_8702_), .Y(_8640_) );
	NAND3X1 NAND3X1_466 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .B(scheduler_block_scheduler_ctr_1_bF_buf2), .C(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_2_), .Y(_8641_) );
	NAND3X1 NAND3X1_467 ( .A(_8641_), .B(_8639_), .C(_8640_), .Y(_8642_) );
	NAND2X1 NAND2X1_1833 ( .A(_8701__bF_buf1), .B(_8642_), .Y(_8643_) );
	NAND2X1 NAND2X1_1834 ( .A(_8638_), .B(_8643_), .Y(_8610__6_) );
	OAI21X1 OAI21X1_308 ( .A(_8699_), .B(rst_bF_buf3), .C(input_selector_block_input_selector_i_3__input_selector_j_1__input_selector_r_3_), .Y(_8644_) );
	NAND3X1 NAND3X1_468 ( .A(scheduler_block_scheduler_ctr_1_bF_buf1), .B(input_selector_block_input_selector_i_1__input_selector_j_1__input_selector_r_3_), .C(_8705_), .Y(_8645_) );
	NAND3X1 NAND3X1_469 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(input_selector_block_input_selector_i_2__input_selector_j_1__input_selector_r_3_), .C(_8702_), .Y(_8646_) );
	NAND3X1 NAND3X1_470 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf0), .C(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_3_), .Y(_8647_) );
	NAND3X1 NAND3X1_471 ( .A(_8647_), .B(_8645_), .C(_8646_), .Y(_8648_) );
	NAND2X1 NAND2X1_1835 ( .A(_8701__bF_buf0), .B(_8648_), .Y(_8649_) );
	NAND2X1 NAND2X1_1836 ( .A(_8644_), .B(_8649_), .Y(_8610__7_) );
	OAI21X1 OAI21X1_309 ( .A(_8699_), .B(rst_bF_buf2), .C(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_0_), .Y(_8650_) );
	NAND3X1 NAND3X1_472 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_0_), .C(_8702_), .Y(_8651_) );
	NAND3X1 NAND3X1_473 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(scheduler_block_scheduler_ctr_1_bF_buf5), .C(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_0_), .Y(_8652_) );
	NAND3X1 NAND3X1_474 ( .A(scheduler_block_scheduler_ctr_1_bF_buf4), .B(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_0_), .C(_8705_), .Y(_8653_) );
	NAND3X1 NAND3X1_475 ( .A(_8652_), .B(_8651_), .C(_8653_), .Y(_8654_) );
	NAND2X1 NAND2X1_1837 ( .A(_8701__bF_buf3), .B(_8654_), .Y(_8655_) );
	NAND2X1 NAND2X1_1838 ( .A(_8650_), .B(_8655_), .Y(_8610__8_) );
	OAI21X1 OAI21X1_310 ( .A(_8699_), .B(rst_bF_buf1), .C(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_1_), .Y(_8656_) );
	NAND3X1 NAND3X1_476 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_1_), .C(_8702_), .Y(_8657_) );
	NAND3X1 NAND3X1_477 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .B(scheduler_block_scheduler_ctr_1_bF_buf3), .C(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_1_), .Y(_8658_) );
	NAND3X1 NAND3X1_478 ( .A(scheduler_block_scheduler_ctr_1_bF_buf2), .B(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_1_), .C(_8705_), .Y(_8659_) );
	NAND3X1 NAND3X1_479 ( .A(_8658_), .B(_8657_), .C(_8659_), .Y(_8660_) );
	NAND2X1 NAND2X1_1839 ( .A(_8701__bF_buf2), .B(_8660_), .Y(_8661_) );
	NAND2X1 NAND2X1_1840 ( .A(_8656_), .B(_8661_), .Y(_8610__9_) );
	OAI21X1 OAI21X1_311 ( .A(_8699_), .B(rst_bF_buf0), .C(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_2_), .Y(_8662_) );
	NAND3X1 NAND3X1_480 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_2_), .C(_8702_), .Y(_8663_) );
	NAND3X1 NAND3X1_481 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf1), .C(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_2_), .Y(_8664_) );
	NAND3X1 NAND3X1_482 ( .A(scheduler_block_scheduler_ctr_1_bF_buf0), .B(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_2_), .C(_8705_), .Y(_8665_) );
	NAND3X1 NAND3X1_483 ( .A(_8664_), .B(_8663_), .C(_8665_), .Y(_8666_) );
	NAND2X1 NAND2X1_1841 ( .A(_8701__bF_buf1), .B(_8666_), .Y(_8667_) );
	NAND2X1 NAND2X1_1842 ( .A(_8662_), .B(_8667_), .Y(_8610__10_) );
	OAI21X1 OAI21X1_312 ( .A(_8699_), .B(rst_bF_buf3), .C(input_selector_block_input_selector_i_3__input_selector_j_2__input_selector_r_3_), .Y(_8668_) );
	NAND3X1 NAND3X1_484 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(input_selector_block_input_selector_i_2__input_selector_j_2__input_selector_r_3_), .C(_8702_), .Y(_8669_) );
	NAND3X1 NAND3X1_485 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(scheduler_block_scheduler_ctr_1_bF_buf5), .C(input_selector_block_input_selector_i_0__input_selector_j_2__input_selector_r_3_), .Y(_8670_) );
	NAND3X1 NAND3X1_486 ( .A(scheduler_block_scheduler_ctr_1_bF_buf4), .B(input_selector_block_input_selector_i_1__input_selector_j_2__input_selector_r_3_), .C(_8705_), .Y(_8671_) );
	NAND3X1 NAND3X1_487 ( .A(_8670_), .B(_8669_), .C(_8671_), .Y(_8672_) );
	NAND2X1 NAND2X1_1843 ( .A(_8701__bF_buf0), .B(_8672_), .Y(_8673_) );
	NAND2X1 NAND2X1_1844 ( .A(_8668_), .B(_8673_), .Y(_8610__11_) );
	OAI21X1 OAI21X1_313 ( .A(_8699_), .B(rst_bF_buf2), .C(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_0_), .Y(_8674_) );
	NAND3X1 NAND3X1_488 ( .A(scheduler_block_scheduler_ctr_1_bF_buf3), .B(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_0_), .C(_8705_), .Y(_8675_) );
	NAND3X1 NAND3X1_489 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_0_), .C(_8702_), .Y(_8676_) );
	NAND3X1 NAND3X1_490 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .B(scheduler_block_scheduler_ctr_1_bF_buf2), .C(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_0_), .Y(_8677_) );
	NAND3X1 NAND3X1_491 ( .A(_8677_), .B(_8675_), .C(_8676_), .Y(_8678_) );
	NAND2X1 NAND2X1_1845 ( .A(_8701__bF_buf3), .B(_8678_), .Y(_8679_) );
	NAND2X1 NAND2X1_1846 ( .A(_8674_), .B(_8679_), .Y(_8610__12_) );
	OAI21X1 OAI21X1_314 ( .A(_8699_), .B(rst_bF_buf1), .C(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_1_), .Y(_8680_) );
	NAND3X1 NAND3X1_492 ( .A(scheduler_block_scheduler_ctr_1_bF_buf1), .B(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_1_), .C(_8705_), .Y(_8681_) );
	NAND3X1 NAND3X1_493 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_1_), .C(_8702_), .Y(_8682_) );
	NAND3X1 NAND3X1_494 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf0), .C(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_1_), .Y(_8683_) );
	NAND3X1 NAND3X1_495 ( .A(_8683_), .B(_8681_), .C(_8682_), .Y(_8684_) );
	NAND2X1 NAND2X1_1847 ( .A(_8701__bF_buf2), .B(_8684_), .Y(_8685_) );
	NAND2X1 NAND2X1_1848 ( .A(_8680_), .B(_8685_), .Y(_8610__13_) );
	OAI21X1 OAI21X1_315 ( .A(_8699_), .B(rst_bF_buf0), .C(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_2_), .Y(_8686_) );
	NAND3X1 NAND3X1_496 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_2_), .C(_8702_), .Y(_8687_) );
	NAND3X1 NAND3X1_497 ( .A(scheduler_block_scheduler_ctr_0_bF_buf4), .B(scheduler_block_scheduler_ctr_1_bF_buf5), .C(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_2_), .Y(_8688_) );
	NAND3X1 NAND3X1_498 ( .A(scheduler_block_scheduler_ctr_1_bF_buf4), .B(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_2_), .C(_8705_), .Y(_8689_) );
	NAND3X1 NAND3X1_499 ( .A(_8688_), .B(_8687_), .C(_8689_), .Y(_8690_) );
	NAND2X1 NAND2X1_1849 ( .A(_8701__bF_buf1), .B(_8690_), .Y(_8691_) );
	NAND2X1 NAND2X1_1850 ( .A(_8686_), .B(_8691_), .Y(_8610__14_) );
	OAI21X1 OAI21X1_316 ( .A(_8699_), .B(rst_bF_buf3), .C(input_selector_block_input_selector_i_3__input_selector_j_3__input_selector_r_3_), .Y(_8692_) );
	NAND3X1 NAND3X1_500 ( .A(scheduler_block_scheduler_ctr_1_bF_buf3), .B(input_selector_block_input_selector_i_1__input_selector_j_3__input_selector_r_3_), .C(_8705_), .Y(_8693_) );
	NAND3X1 NAND3X1_501 ( .A(scheduler_block_scheduler_ctr_0_bF_buf3), .B(input_selector_block_input_selector_i_2__input_selector_j_3__input_selector_r_3_), .C(_8702_), .Y(_8694_) );
	NAND3X1 NAND3X1_502 ( .A(scheduler_block_scheduler_ctr_0_bF_buf2), .B(scheduler_block_scheduler_ctr_1_bF_buf2), .C(input_selector_block_input_selector_i_0__input_selector_j_3__input_selector_r_3_), .Y(_8695_) );
	NAND3X1 NAND3X1_503 ( .A(_8695_), .B(_8693_), .C(_8694_), .Y(_8696_) );
	NAND2X1 NAND2X1_1851 ( .A(_8701__bF_buf0), .B(_8696_), .Y(_8697_) );
	NAND2X1 NAND2X1_1852 ( .A(_8692_), .B(_8697_), .Y(_8610__15_) );
	NOR2X1 NOR2X1_1047 ( .A(scheduler_block_scheduler_ctr_0_bF_buf1), .B(rst_bF_buf2), .Y(_8609__0_) );
	OAI21X1 OAI21X1_317 ( .A(scheduler_block_scheduler_ctr_0_bF_buf0), .B(scheduler_block_scheduler_ctr_1_bF_buf1), .C(_8701__bF_buf3), .Y(_8698_) );
	AOI21X1 AOI21X1_214 ( .A(scheduler_block_scheduler_ctr_0_bF_buf5), .B(scheduler_block_scheduler_ctr_1_bF_buf0), .C(_8698_), .Y(_8609__1_) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf42), .D(_8610__0_), .Q(scheduler_block_data_out_0_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf41), .D(_8610__1_), .Q(scheduler_block_data_out_1_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf40), .D(_8610__2_), .Q(scheduler_block_data_out_2_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf39), .D(_8610__3_), .Q(scheduler_block_data_out_3_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf38), .D(_8610__4_), .Q(scheduler_block_data_out_4_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf37), .D(_8610__5_), .Q(scheduler_block_data_out_5_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf36), .D(_8610__6_), .Q(scheduler_block_data_out_6_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf35), .D(_8610__7_), .Q(scheduler_block_data_out_7_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf34), .D(_8610__8_), .Q(scheduler_block_data_out_8_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf33), .D(_8610__9_), .Q(scheduler_block_data_out_9_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf32), .D(_8610__10_), .Q(scheduler_block_data_out_10_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf31), .D(_8610__11_), .Q(scheduler_block_data_out_11_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf30), .D(_8610__12_), .Q(scheduler_block_data_out_12_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf29), .D(_8610__13_), .Q(scheduler_block_data_out_13_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf28), .D(_8610__14_), .Q(scheduler_block_data_out_14_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf27), .D(_8610__15_), .Q(scheduler_block_data_out_15_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf26), .D(_8609__0_), .Q(scheduler_block_scheduler_ctr_0_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf25), .D(_8609__1_), .Q(scheduler_block_scheduler_ctr_1_) );
	BUFX2 BUFX2_32 ( .A(_0__0_), .Y(data_out[0]) );
	BUFX2 BUFX2_33 ( .A(_0__1_), .Y(data_out[1]) );
	BUFX2 BUFX2_34 ( .A(_0__2_), .Y(data_out[2]) );
	BUFX2 BUFX2_35 ( .A(_0__3_), .Y(data_out[3]) );
	BUFX2 BUFX2_36 ( .A(_0__4_), .Y(data_out[4]) );
	BUFX2 BUFX2_37 ( .A(_0__5_), .Y(data_out[5]) );
	BUFX2 BUFX2_38 ( .A(_0__6_), .Y(data_out[6]) );
	BUFX2 BUFX2_39 ( .A(_0__7_), .Y(data_out[7]) );
	BUFX2 BUFX2_40 ( .A(_0__8_), .Y(data_out[8]) );
	BUFX2 BUFX2_41 ( .A(_0__9_), .Y(data_out[9]) );
	BUFX2 BUFX2_42 ( .A(_0__10_), .Y(data_out[10]) );
	BUFX2 BUFX2_43 ( .A(_0__11_), .Y(data_out[11]) );
	BUFX2 BUFX2_44 ( .A(_0__12_), .Y(data_out[12]) );
	BUFX2 BUFX2_45 ( .A(_0__13_), .Y(data_out[13]) );
	BUFX2 BUFX2_46 ( .A(_0__14_), .Y(data_out[14]) );
	BUFX2 BUFX2_47 ( .A(_0__15_), .Y(data_out[15]) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf24), .D(wRegs0[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf23), .D(wRegs0[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf22), .D(wRegs0[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf21), .D(wRegs0[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf20), .D(wRegs0[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf19), .D(wRegs0[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf18), .D(wRegs0[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf17), .D(wRegs0[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf16), .D(wRegs0[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf15), .D(wRegs0[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf14), .D(wRegs0[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf13), .D(wRegs0[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf12), .D(wRegs0[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf11), .D(wRegs0[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf10), .D(wRegs0[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf9), .D(wRegs0[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf8), .D(wRegs0[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf7), .D(wRegs0[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf6), .D(wRegs0[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf5), .D(wRegs0[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf4), .D(wRegs0[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf3), .D(wRegs0[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf2), .D(wRegs0[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf1), .D(wRegs0[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf0), .D(wRegs0[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf42), .D(wRegs0[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf41), .D(wRegs0[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf40), .D(wRegs0[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf39), .D(wRegs0[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf38), .D(wRegs0[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf37), .D(wRegs0[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf36), .D(wRegs0[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf35), .D(wRegs1[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf34), .D(wRegs1[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf33), .D(wRegs1[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf32), .D(wRegs1[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf31), .D(wRegs1[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf30), .D(wRegs1[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf29), .D(wRegs1[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf28), .D(wRegs1[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf27), .D(wRegs1[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf26), .D(wRegs1[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf25), .D(wRegs1[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf24), .D(wRegs1[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf23), .D(wRegs1[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf22), .D(wRegs1[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf21), .D(wRegs1[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf20), .D(wRegs1[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf19), .D(wRegs1[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf18), .D(wRegs1[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf17), .D(wRegs1[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf16), .D(wRegs1[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf15), .D(wRegs1[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf14), .D(wRegs1[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf13), .D(wRegs1[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf12), .D(wRegs1[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf11), .D(wRegs1[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf10), .D(wRegs1[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf9), .D(wRegs1[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf8), .D(wRegs1[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf7), .D(wRegs1[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf6), .D(wRegs1[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_) );
	DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf5), .D(wRegs1[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_) );
	DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf4), .D(wRegs1[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_) );
	DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf3), .D(wRegs2[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_) );
	DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf2), .D(wRegs2[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_) );
	DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf1), .D(wRegs2[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_) );
	DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf0), .D(wRegs2[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_) );
	DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf42), .D(wRegs2[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_) );
	DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf41), .D(wRegs2[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_) );
	DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf40), .D(wRegs2[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_) );
	DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf39), .D(wRegs2[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_) );
	DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf38), .D(wRegs2[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_) );
	DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf37), .D(wRegs2[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_) );
	DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf36), .D(wRegs2[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_) );
	DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf35), .D(wRegs2[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_) );
	DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf34), .D(wRegs2[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_) );
	DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf33), .D(wRegs2[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_) );
	DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf32), .D(wRegs2[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_) );
	DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf31), .D(wRegs2[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_) );
	DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf30), .D(wRegs2[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_) );
	DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf29), .D(wRegs2[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_) );
	DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf28), .D(wRegs2[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_) );
	DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf27), .D(wRegs2[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_) );
	DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf26), .D(wRegs2[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_) );
	DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf25), .D(wRegs2[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_) );
	DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf24), .D(wRegs2[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_) );
	DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf23), .D(wRegs2[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_) );
	DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf22), .D(wRegs2[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_) );
	DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf21), .D(wRegs2[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_) );
	DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf20), .D(wRegs2[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_) );
	DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf19), .D(wRegs2[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_) );
	DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf18), .D(wRegs2[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_) );
	DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf17), .D(wRegs2[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_) );
	DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf16), .D(wRegs2[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_) );
	DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf15), .D(wRegs2[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_) );
	DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf14), .D(wRegs3[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_) );
	DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf13), .D(wRegs3[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_) );
	DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf12), .D(wRegs3[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_) );
	DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf11), .D(wRegs3[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_) );
	DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf10), .D(wRegs3[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_) );
	DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf9), .D(wRegs3[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_) );
	DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf8), .D(wRegs3[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_) );
	DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf7), .D(wRegs3[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_) );
	DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf6), .D(wRegs3[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_) );
	DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf5), .D(wRegs3[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_) );
	DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf4), .D(wRegs3[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_) );
	DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf3), .D(wRegs3[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_) );
	DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf2), .D(wRegs3[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_) );
	DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf1), .D(wRegs3[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_) );
	DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf0), .D(wRegs3[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_) );
	DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf42), .D(wRegs3[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_) );
	DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf41), .D(wRegs3[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_) );
	DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf40), .D(wRegs3[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_) );
	DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf39), .D(wRegs3[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_) );
	DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf38), .D(wRegs3[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_) );
	DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf37), .D(wRegs3[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_) );
	DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf36), .D(wRegs3[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_) );
	DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf35), .D(wRegs3[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_) );
	DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf34), .D(wRegs3[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_) );
	DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf33), .D(wRegs3[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_) );
	DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf32), .D(wRegs3[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_) );
	DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf31), .D(wRegs3[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_) );
	DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf30), .D(wRegs3[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_) );
	DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf29), .D(wRegs3[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_) );
	DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf28), .D(wRegs3[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_) );
	DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf27), .D(wRegs3[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_) );
	DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf26), .D(wRegs3[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_) );
	DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf25), .D(wRegs4[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_) );
	DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf24), .D(wRegs4[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_) );
	DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf23), .D(wRegs4[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_) );
	DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf22), .D(wRegs4[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_) );
	DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf21), .D(wRegs4[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_) );
	DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf20), .D(wRegs4[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_) );
	DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf19), .D(wRegs4[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_) );
	DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf18), .D(wRegs4[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_) );
	DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf17), .D(wRegs4[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_) );
	DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf16), .D(wRegs4[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_) );
	DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf15), .D(wRegs4[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_) );
	DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf14), .D(wRegs4[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_) );
	DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf13), .D(wRegs4[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_) );
	DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf12), .D(wRegs4[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_) );
	DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf11), .D(wRegs4[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_) );
	DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf10), .D(wRegs4[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_) );
	DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf9), .D(wRegs4[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_) );
	DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf8), .D(wRegs4[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_) );
	DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf7), .D(wRegs4[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_) );
	DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf6), .D(wRegs4[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_) );
	DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf5), .D(wRegs4[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_) );
	DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf4), .D(wRegs4[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_) );
	DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf3), .D(wRegs4[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_) );
	DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf2), .D(wRegs4[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_) );
	DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf1), .D(wRegs4[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_) );
	DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf0), .D(wRegs4[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_) );
	DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf42), .D(wRegs4[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_) );
	DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf41), .D(wRegs4[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_) );
	DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf40), .D(wRegs4[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_) );
	DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf39), .D(wRegs4[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_) );
	DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf38), .D(wRegs4[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_) );
	DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf37), .D(wRegs4[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_) );
	DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf36), .D(wRegs5[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_) );
	DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf35), .D(wRegs5[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_) );
	DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf34), .D(wRegs5[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_) );
	DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf33), .D(wRegs5[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_) );
	DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf32), .D(wRegs5[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_) );
	DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf31), .D(wRegs5[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_) );
	DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf30), .D(wRegs5[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_) );
	DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf29), .D(wRegs5[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_) );
	DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf28), .D(wRegs5[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_) );
	DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf27), .D(wRegs5[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_) );
	DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf26), .D(wRegs5[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_) );
	DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf25), .D(wRegs5[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_) );
	DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf24), .D(wRegs5[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_) );
	DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf23), .D(wRegs5[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_) );
	DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf22), .D(wRegs5[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_) );
	DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf21), .D(wRegs5[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_) );
	DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf20), .D(wRegs5[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_) );
	DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf19), .D(wRegs5[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_) );
	DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf18), .D(wRegs5[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_) );
	DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf17), .D(wRegs5[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_) );
	DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf16), .D(wRegs5[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_) );
	DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf15), .D(wRegs5[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_) );
	DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf14), .D(wRegs5[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_) );
	DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf13), .D(wRegs5[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_) );
	DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf12), .D(wRegs5[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_) );
	DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf11), .D(wRegs5[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_) );
	DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf10), .D(wRegs5[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_) );
	DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf9), .D(wRegs5[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_) );
	DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf8), .D(wRegs5[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_) );
	DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf7), .D(wRegs5[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_) );
	DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf6), .D(wRegs5[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_) );
	DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf5), .D(wRegs5[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_) );
	DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf4), .D(wRegs6[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_) );
	DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf3), .D(wRegs6[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_) );
	DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf2), .D(wRegs6[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_) );
	DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf1), .D(wRegs6[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_) );
	DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf0), .D(wRegs6[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_) );
	DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf42), .D(wRegs6[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_) );
	DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf41), .D(wRegs6[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_) );
	DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf40), .D(wRegs6[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_) );
	DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf39), .D(wRegs6[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_) );
	DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf38), .D(wRegs6[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_) );
	DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf37), .D(wRegs6[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_) );
	DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf36), .D(wRegs6[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_) );
	DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf35), .D(wRegs6[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_) );
	DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf34), .D(wRegs6[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_) );
	DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf33), .D(wRegs6[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_) );
	DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf32), .D(wRegs6[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_) );
	DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf31), .D(wRegs6[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_) );
	DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf30), .D(wRegs6[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_) );
	DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf29), .D(wRegs6[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_) );
	DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf28), .D(wRegs6[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_) );
	DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf27), .D(wRegs6[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_) );
	DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf26), .D(wRegs6[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_) );
	DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf25), .D(wRegs6[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_) );
	DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf24), .D(wRegs6[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_) );
	DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf23), .D(wRegs6[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_) );
	DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf22), .D(wRegs6[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_) );
	DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf21), .D(wRegs6[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_) );
	DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf20), .D(wRegs6[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_) );
	DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf19), .D(wRegs6[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_) );
	DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf18), .D(wRegs6[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_) );
	DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf17), .D(wRegs6[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_) );
	DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf16), .D(wRegs6[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_) );
	DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf15), .D(wRegs7[0]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_) );
	DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf14), .D(wRegs7[1]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_) );
	DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf13), .D(wRegs7[2]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_) );
	DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf12), .D(wRegs7[3]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_) );
	DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf11), .D(wRegs7[4]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_) );
	DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf10), .D(wRegs7[5]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_) );
	DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf9), .D(wRegs7[6]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_) );
	DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf8), .D(wRegs7[7]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_) );
	DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf7), .D(wRegs7[8]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_) );
	DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf6), .D(wRegs7[9]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_) );
	DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf5), .D(wRegs7[10]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_) );
	DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf4), .D(wRegs7[11]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_) );
	DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf3), .D(wRegs7[12]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_) );
	DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf2), .D(wRegs7[13]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_) );
	DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf1), .D(wRegs7[14]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_) );
	DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf0), .D(wRegs7[15]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_) );
	DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf42), .D(wRegs7[16]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_) );
	DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf41), .D(wRegs7[17]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_) );
	DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf40), .D(wRegs7[18]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_) );
	DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf39), .D(wRegs7[19]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_) );
	DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf38), .D(wRegs7[20]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_) );
	DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf37), .D(wRegs7[21]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_) );
	DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf36), .D(wRegs7[22]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_) );
	DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf35), .D(wRegs7[23]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_) );
	DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf34), .D(wRegs7[24]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_) );
	DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf33), .D(wRegs7[25]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_) );
	DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf32), .D(wRegs7[26]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_) );
	DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf31), .D(wRegs7[27]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_) );
	DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf30), .D(wRegs7[28]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_) );
	DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf29), .D(wRegs7[29]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_) );
	DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf28), .D(wRegs7[30]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_) );
	DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf27), .D(wRegs7[31]), .Q(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_) );
	DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf26), .D(scheduler_block_data_out_0_), .Q(_0__0_) );
	DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf25), .D(scheduler_block_data_out_1_), .Q(_0__1_) );
	DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf24), .D(scheduler_block_data_out_2_), .Q(_0__2_) );
	DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf23), .D(scheduler_block_data_out_3_), .Q(_0__3_) );
	DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf22), .D(scheduler_block_data_out_4_), .Q(_0__4_) );
	DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf21), .D(scheduler_block_data_out_5_), .Q(_0__5_) );
	DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf20), .D(scheduler_block_data_out_6_), .Q(_0__6_) );
	DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf19), .D(scheduler_block_data_out_7_), .Q(_0__7_) );
	DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf18), .D(scheduler_block_data_out_8_), .Q(_0__8_) );
	DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf17), .D(scheduler_block_data_out_9_), .Q(_0__9_) );
	DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf16), .D(scheduler_block_data_out_10_), .Q(_0__10_) );
	DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf15), .D(scheduler_block_data_out_11_), .Q(_0__11_) );
	DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf14), .D(scheduler_block_data_out_12_), .Q(_0__12_) );
	DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf13), .D(scheduler_block_data_out_13_), .Q(_0__13_) );
	DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf12), .D(scheduler_block_data_out_14_), .Q(_0__14_) );
	DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf11), .D(scheduler_block_data_out_15_), .Q(_0__15_) );
	INVX1 INVX1_1130 ( .A(wSelec[0]), .Y(_1_) );
	NOR2X1 NOR2X1_1048 ( .A(wBusy_bF_buf0), .B(_1_), .Y(_2_) );
	INVX1 INVX1_1131 ( .A(_2_), .Y(_3_) );
	INVX1 INVX1_1132 ( .A(wSelec[10]), .Y(_4_) );
	NAND2X1 NAND2X1_1853 ( .A(wSelec[9]), .B(_4_), .Y(_5_) );
	INVX2 INVX2_29 ( .A(_5_), .Y(_6_) );
	OR2X2 OR2X2_100 ( .A(wSelec[6]), .B(wSelec[5]), .Y(_7_) );
	INVX1 INVX1_1133 ( .A(wSelec[8]), .Y(_8_) );
	NAND2X1 NAND2X1_1854 ( .A(wSelec[7]), .B(_8_), .Y(_9_) );
	NOR2X1 NOR2X1_1049 ( .A(_7_), .B(_9_), .Y(_10_) );
	AND2X2 AND2X2_198 ( .A(_10_), .B(_6_), .Y(_11_) );
	AOI21X1 AOI21X1_215 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_11_), .C(_3_), .Y(_12_) );
	INVX1 INVX1_1134 ( .A(wSelec[6]), .Y(_13_) );
	NAND2X1 NAND2X1_1855 ( .A(wSelec[5]), .B(_13_), .Y(_14_) );
	OR2X2 OR2X2_101 ( .A(wSelec[7]), .B(wSelec[8]), .Y(_15_) );
	NOR2X1 NOR2X1_1050 ( .A(_15_), .B(_14_), .Y(_16_) );
	NAND2X1 NAND2X1_1856 ( .A(_6_), .B(_16_), .Y(_17_) );
	INVX1 INVX1_1135 ( .A(_17_), .Y(_18_) );
	INVX1 INVX1_1136 ( .A(wSelec[5]), .Y(_19_) );
	NAND2X1 NAND2X1_1857 ( .A(wSelec[6]), .B(_19_), .Y(_20_) );
	INVX1 INVX1_1137 ( .A(wSelec[7]), .Y(_21_) );
	NAND2X1 NAND2X1_1858 ( .A(wSelec[8]), .B(_21_), .Y(_22_) );
	NOR2X1 NOR2X1_1051 ( .A(_20_), .B(_22_), .Y(_23_) );
	NAND2X1 NAND2X1_1859 ( .A(wSelec[9]), .B(wSelec[10]), .Y(_24_) );
	INVX1 INVX1_1138 ( .A(_24_), .Y(_25_) );
	NAND2X1 NAND2X1_1860 ( .A(_25_), .B(_23_), .Y(_26_) );
	INVX1 INVX1_1139 ( .A(_26_), .Y(_27_) );
	AOI22X1 AOI22X1_1419 ( .A(_18_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_27_), .Y(_28_) );
	OR2X2 OR2X2_102 ( .A(_14_), .B(_15_), .Y(_29_) );
	OR2X2 OR2X2_103 ( .A(wSelec[9]), .B(wSelec[10]), .Y(_30_) );
	NOR2X1 NOR2X1_1052 ( .A(_30_), .B(_29_), .Y(_31_) );
	NOR2X1 NOR2X1_1053 ( .A(_9_), .B(_14_), .Y(_32_) );
	INVX1 INVX1_1140 ( .A(wSelec[9]), .Y(_33_) );
	NAND2X1 NAND2X1_1861 ( .A(wSelec[10]), .B(_33_), .Y(_34_) );
	INVX2 INVX2_30 ( .A(_34_), .Y(_35_) );
	NAND2X1 NAND2X1_1862 ( .A(_35_), .B(_32_), .Y(_36_) );
	INVX1 INVX1_1141 ( .A(_36_), .Y(_37_) );
	AOI22X1 AOI22X1_1420 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_31_), .C(_37_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_38_) );
	NAND3X1 NAND3X1_504 ( .A(_12_), .B(_38_), .C(_28_), .Y(_39_) );
	NOR2X1 NOR2X1_1054 ( .A(wSelec[6]), .B(wSelec[5]), .Y(_40_) );
	NOR2X1 NOR2X1_1055 ( .A(wSelec[7]), .B(wSelec[8]), .Y(_41_) );
	NAND2X1 NAND2X1_1863 ( .A(_40_), .B(_41_), .Y(_42_) );
	NOR2X1 NOR2X1_1056 ( .A(_5_), .B(_42_), .Y(_43_) );
	NAND2X1 NAND2X1_1864 ( .A(wSelec[6]), .B(wSelec[5]), .Y(_44_) );
	NOR3X1 NOR3X1_745 ( .A(_15_), .B(_44_), .C(_5_), .Y(_45_) );
	AOI22X1 AOI22X1_1421 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_45_), .C(_43_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_46_) );
	INVX1 INVX1_1142 ( .A(_30_), .Y(_47_) );
	NOR2X1 NOR2X1_1057 ( .A(_15_), .B(_20_), .Y(_48_) );
	AND2X2 AND2X2_199 ( .A(_48_), .B(_47_), .Y(_49_) );
	NAND2X1 NAND2X1_1865 ( .A(wSelec[7]), .B(wSelec[8]), .Y(_50_) );
	NOR3X1 NOR3X1_746 ( .A(_24_), .B(_44_), .C(_50_), .Y(_51_) );
	AOI22X1 AOI22X1_1422 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_51_), .C(_49_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_52_) );
	INVX1 INVX1_1143 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_53_) );
	INVX1 INVX1_1144 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_54_) );
	NOR2X1 NOR2X1_1058 ( .A(_14_), .B(_22_), .Y(_55_) );
	NAND2X1 NAND2X1_1866 ( .A(_25_), .B(_55_), .Y(_56_) );
	NOR2X1 NOR2X1_1059 ( .A(_44_), .B(_50_), .Y(_57_) );
	NAND2X1 NAND2X1_1867 ( .A(_57_), .B(_35_), .Y(_58_) );
	OAI22X1 OAI22X1_241 ( .A(_53_), .B(_58_), .C(_56_), .D(_54_), .Y(_59_) );
	INVX1 INVX1_1145 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_60_) );
	NOR3X1 NOR3X1_747 ( .A(_5_), .B(_20_), .C(_22_), .Y(_61_) );
	NAND2X1 NAND2X1_1868 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_61_), .Y(_62_) );
	NOR2X1 NOR2X1_1060 ( .A(_44_), .B(_9_), .Y(_63_) );
	NAND2X1 NAND2X1_1869 ( .A(_35_), .B(_63_), .Y(_64_) );
	OAI21X1 OAI21X1_318 ( .A(_60_), .B(_64_), .C(_62_), .Y(_65_) );
	NOR2X1 NOR2X1_1061 ( .A(_59_), .B(_65_), .Y(_66_) );
	NAND3X1 NAND3X1_505 ( .A(_46_), .B(_52_), .C(_66_), .Y(_67_) );
	INVX1 INVX1_1146 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_68_) );
	INVX1 INVX1_1147 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_69_) );
	NOR2X1 NOR2X1_1062 ( .A(_9_), .B(_20_), .Y(_70_) );
	NAND2X1 NAND2X1_1870 ( .A(_6_), .B(_70_), .Y(_71_) );
	NOR2X1 NOR2X1_1063 ( .A(_7_), .B(_22_), .Y(_72_) );
	NAND2X1 NAND2X1_1871 ( .A(_6_), .B(_72_), .Y(_73_) );
	OAI22X1 OAI22X1_242 ( .A(_73_), .B(_68_), .C(_69_), .D(_71_), .Y(_74_) );
	INVX1 INVX1_1148 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_75_) );
	INVX1 INVX1_1149 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_76_) );
	NAND2X1 NAND2X1_1872 ( .A(_35_), .B(_70_), .Y(_77_) );
	NOR2X1 NOR2X1_1064 ( .A(_44_), .B(_15_), .Y(_78_) );
	NAND2X1 NAND2X1_1873 ( .A(_35_), .B(_78_), .Y(_79_) );
	OAI22X1 OAI22X1_243 ( .A(_75_), .B(_79_), .C(_77_), .D(_76_), .Y(_80_) );
	NOR2X1 NOR2X1_1065 ( .A(_80_), .B(_74_), .Y(_81_) );
	NOR3X1 NOR3X1_748 ( .A(_14_), .B(_50_), .C(_34_), .Y(_82_) );
	NAND2X1 NAND2X1_1874 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_82_), .Y(_83_) );
	NOR3X1 NOR3X1_749 ( .A(_22_), .B(_44_), .C(_34_), .Y(_84_) );
	NAND2X1 NAND2X1_1875 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_84_), .Y(_85_) );
	NAND2X1 NAND2X1_1876 ( .A(_83_), .B(_85_), .Y(_86_) );
	INVX1 INVX1_1150 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_87_) );
	NAND2X1 NAND2X1_1877 ( .A(_25_), .B(_10_), .Y(_88_) );
	NOR3X1 NOR3X1_750 ( .A(_20_), .B(_22_), .C(_34_), .Y(_89_) );
	NAND2X1 NAND2X1_1878 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_89_), .Y(_90_) );
	OAI21X1 OAI21X1_319 ( .A(_87_), .B(_88_), .C(_90_), .Y(_91_) );
	NOR2X1 NOR2X1_1066 ( .A(_86_), .B(_91_), .Y(_92_) );
	NAND2X1 NAND2X1_1879 ( .A(_81_), .B(_92_), .Y(_93_) );
	NOR3X1 NOR3X1_751 ( .A(_39_), .B(_93_), .C(_67_), .Y(_94_) );
	NAND2X1 NAND2X1_1880 ( .A(_6_), .B(_63_), .Y(_95_) );
	INVX1 INVX1_1151 ( .A(_95_), .Y(_96_) );
	INVX1 INVX1_1152 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_97_) );
	NOR3X1 NOR3X1_752 ( .A(_7_), .B(_30_), .C(_9_), .Y(_98_) );
	NAND2X1 NAND2X1_1881 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_98_), .Y(_99_) );
	NAND2X1 NAND2X1_1882 ( .A(_47_), .B(_70_), .Y(_100_) );
	OAI21X1 OAI21X1_320 ( .A(_100_), .B(_97_), .C(_99_), .Y(_101_) );
	AOI21X1 AOI21X1_216 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_96_), .C(_101_), .Y(_102_) );
	INVX1 INVX1_1153 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_103_) );
	INVX1 INVX1_1154 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_104_) );
	NOR2X1 NOR2X1_1067 ( .A(_50_), .B(_7_), .Y(_105_) );
	NAND2X1 NAND2X1_1883 ( .A(_6_), .B(_105_), .Y(_106_) );
	NAND2X1 NAND2X1_1884 ( .A(_47_), .B(_32_), .Y(_107_) );
	OAI22X1 OAI22X1_244 ( .A(_104_), .B(_106_), .C(_107_), .D(_103_), .Y(_108_) );
	INVX1 INVX1_1155 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_109_) );
	INVX1 INVX1_1156 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_110_) );
	NAND2X1 NAND2X1_1885 ( .A(_6_), .B(_32_), .Y(_111_) );
	NAND2X1 NAND2X1_1886 ( .A(_47_), .B(_78_), .Y(_112_) );
	OAI22X1 OAI22X1_245 ( .A(_109_), .B(_112_), .C(_111_), .D(_110_), .Y(_113_) );
	NOR2X1 NOR2X1_1068 ( .A(_108_), .B(_113_), .Y(_114_) );
	INVX1 INVX1_1157 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_115_) );
	NOR3X1 NOR3X1_753 ( .A(_30_), .B(_44_), .C(_9_), .Y(_116_) );
	NAND2X1 NAND2X1_1887 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_116_), .Y(_117_) );
	OR2X2 OR2X2_104 ( .A(_42_), .B(_24_), .Y(_118_) );
	OAI21X1 OAI21X1_321 ( .A(_115_), .B(_118_), .C(_117_), .Y(_119_) );
	INVX1 INVX1_1158 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_120_) );
	INVX1 INVX1_1159 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_121_) );
	NOR2X1 NOR2X1_1069 ( .A(_50_), .B(_20_), .Y(_122_) );
	NAND2X1 NAND2X1_1888 ( .A(_6_), .B(_122_), .Y(_123_) );
	NAND2X1 NAND2X1_1889 ( .A(_25_), .B(_16_), .Y(_124_) );
	OAI22X1 OAI22X1_246 ( .A(_123_), .B(_121_), .C(_120_), .D(_124_), .Y(_125_) );
	NOR2X1 NOR2X1_1070 ( .A(_119_), .B(_125_), .Y(_126_) );
	NAND3X1 NAND3X1_506 ( .A(_102_), .B(_126_), .C(_114_), .Y(_127_) );
	NOR3X1 NOR3X1_754 ( .A(_7_), .B(_15_), .C(_30_), .Y(_128_) );
	NOR3X1 NOR3X1_755 ( .A(_24_), .B(_50_), .C(_14_), .Y(_129_) );
	AOI22X1 AOI22X1_1423 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_128_), .C(_129_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_130_) );
	NOR3X1 NOR3X1_756 ( .A(_24_), .B(_50_), .C(_20_), .Y(_131_) );
	NOR3X1 NOR3X1_757 ( .A(_24_), .B(_44_), .C(_22_), .Y(_132_) );
	AOI22X1 AOI22X1_1424 ( .A(_131_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_132_), .Y(_133_) );
	NAND2X1 NAND2X1_1890 ( .A(_130_), .B(_133_), .Y(_134_) );
	NOR3X1 NOR3X1_758 ( .A(_22_), .B(_7_), .C(_34_), .Y(_135_) );
	NOR3X1 NOR3X1_759 ( .A(_14_), .B(_22_), .C(_34_), .Y(_136_) );
	AOI22X1 AOI22X1_1425 ( .A(_135_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_136_), .Y(_137_) );
	NOR3X1 NOR3X1_760 ( .A(_5_), .B(_50_), .C(_14_), .Y(_138_) );
	NOR3X1 NOR3X1_761 ( .A(_44_), .B(_50_), .C(_5_), .Y(_139_) );
	AOI22X1 AOI22X1_1426 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_139_), .C(_138_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_140_) );
	NAND2X1 NAND2X1_1891 ( .A(_140_), .B(_137_), .Y(_141_) );
	NOR2X1 NOR2X1_1071 ( .A(_134_), .B(_141_), .Y(_142_) );
	NOR3X1 NOR3X1_762 ( .A(_30_), .B(_50_), .C(_14_), .Y(_143_) );
	NOR3X1 NOR3X1_763 ( .A(_30_), .B(_50_), .C(_20_), .Y(_144_) );
	AOI22X1 AOI22X1_1427 ( .A(_143_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_144_), .Y(_145_) );
	NOR3X1 NOR3X1_764 ( .A(_30_), .B(_44_), .C(_22_), .Y(_146_) );
	NOR3X1 NOR3X1_765 ( .A(_5_), .B(_15_), .C(_20_), .Y(_147_) );
	AOI22X1 AOI22X1_1428 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_146_), .C(_147_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_148_) );
	NAND2X1 NAND2X1_1892 ( .A(_145_), .B(_148_), .Y(_149_) );
	NOR3X1 NOR3X1_766 ( .A(_44_), .B(_50_), .C(_30_), .Y(_150_) );
	NOR3X1 NOR3X1_767 ( .A(_20_), .B(_15_), .C(_34_), .Y(_151_) );
	AOI22X1 AOI22X1_1429 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_150_), .C(_151_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_152_) );
	NOR3X1 NOR3X1_768 ( .A(_7_), .B(_15_), .C(_34_), .Y(_153_) );
	NOR3X1 NOR3X1_769 ( .A(_7_), .B(_50_), .C(_34_), .Y(_154_) );
	AOI22X1 AOI22X1_1430 ( .A(_153_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_154_), .Y(_155_) );
	NAND2X1 NAND2X1_1893 ( .A(_155_), .B(_152_), .Y(_156_) );
	NOR2X1 NOR2X1_1072 ( .A(_149_), .B(_156_), .Y(_157_) );
	NAND2X1 NAND2X1_1894 ( .A(_157_), .B(_142_), .Y(_158_) );
	NOR3X1 NOR3X1_770 ( .A(_5_), .B(_44_), .C(_22_), .Y(_159_) );
	NOR3X1 NOR3X1_771 ( .A(_15_), .B(_24_), .C(_20_), .Y(_160_) );
	AOI22X1 AOI22X1_1431 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_160_), .C(_159_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_161_) );
	NOR3X1 NOR3X1_772 ( .A(_9_), .B(_7_), .C(_34_), .Y(_162_) );
	NOR3X1 NOR3X1_773 ( .A(_20_), .B(_50_), .C(_34_), .Y(_163_) );
	AOI22X1 AOI22X1_1432 ( .A(_162_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_163_), .Y(_164_) );
	NAND2X1 NAND2X1_1895 ( .A(_161_), .B(_164_), .Y(_165_) );
	NOR3X1 NOR3X1_774 ( .A(_5_), .B(_14_), .C(_22_), .Y(_166_) );
	NAND2X1 NAND2X1_1896 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_166_), .Y(_167_) );
	NOR3X1 NOR3X1_775 ( .A(_24_), .B(_44_), .C(_9_), .Y(_168_) );
	NAND2X1 NAND2X1_1897 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_168_), .Y(_169_) );
	NOR3X1 NOR3X1_776 ( .A(_7_), .B(_50_), .C(_30_), .Y(_170_) );
	NOR3X1 NOR3X1_777 ( .A(_7_), .B(_24_), .C(_22_), .Y(_171_) );
	AOI22X1 AOI22X1_1433 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_170_), .C(_171_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_172_) );
	NAND3X1 NAND3X1_507 ( .A(_167_), .B(_169_), .C(_172_), .Y(_173_) );
	NOR2X1 NOR2X1_1073 ( .A(_173_), .B(_165_), .Y(_174_) );
	NOR3X1 NOR3X1_778 ( .A(_7_), .B(_30_), .C(_22_), .Y(_175_) );
	NOR3X1 NOR3X1_779 ( .A(_9_), .B(_24_), .C(_14_), .Y(_176_) );
	AOI22X1 AOI22X1_1434 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_175_), .C(_176_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_177_) );
	NOR3X1 NOR3X1_780 ( .A(_9_), .B(_24_), .C(_20_), .Y(_178_) );
	NAND2X1 NAND2X1_1898 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_178_), .Y(_179_) );
	NOR3X1 NOR3X1_781 ( .A(_14_), .B(_15_), .C(_34_), .Y(_180_) );
	NAND2X1 NAND2X1_1899 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_180_), .Y(_181_) );
	NAND3X1 NAND3X1_508 ( .A(_179_), .B(_181_), .C(_177_), .Y(_182_) );
	NOR3X1 NOR3X1_782 ( .A(_14_), .B(_30_), .C(_22_), .Y(_183_) );
	NOR3X1 NOR3X1_783 ( .A(_24_), .B(_50_), .C(_7_), .Y(_184_) );
	AOI22X1 AOI22X1_1435 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_184_), .C(_183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_185_) );
	NOR3X1 NOR3X1_784 ( .A(_20_), .B(_30_), .C(_22_), .Y(_186_) );
	NOR3X1 NOR3X1_785 ( .A(_24_), .B(_44_), .C(_15_), .Y(_187_) );
	AOI22X1 AOI22X1_1436 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_187_), .C(_186_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_188_) );
	NAND2X1 NAND2X1_1900 ( .A(_185_), .B(_188_), .Y(_189_) );
	NOR2X1 NOR2X1_1074 ( .A(_189_), .B(_182_), .Y(_190_) );
	NAND2X1 NAND2X1_1901 ( .A(_174_), .B(_190_), .Y(_191_) );
	NOR3X1 NOR3X1_786 ( .A(_158_), .B(_127_), .C(_191_), .Y(_192_) );
	INVX1 INVX1_1160 ( .A(wSelec[2]), .Y(_193_) );
	NAND2X1 NAND2X1_1902 ( .A(wSelec[1]), .B(_193_), .Y(_194_) );
	INVX1 INVX1_1161 ( .A(wSelec[4]), .Y(_195_) );
	NAND2X1 NAND2X1_1903 ( .A(wSelec[3]), .B(_195_), .Y(_196_) );
	NOR2X1 NOR2X1_1075 ( .A(_194_), .B(_196_), .Y(_197_) );
	NOR2X1 NOR2X1_1076 ( .A(wSelec[2]), .B(wSelec[1]), .Y(_198_) );
	INVX1 INVX1_1162 ( .A(_198_), .Y(_199_) );
	NOR2X1 NOR2X1_1077 ( .A(_196_), .B(_199_), .Y(_200_) );
	AOI22X1 AOI22X1_1437 ( .A(wData[20]), .B(_197_), .C(_200_), .D(wData[16]), .Y(_201_) );
	INVX1 INVX1_1163 ( .A(wSelec[1]), .Y(_202_) );
	NAND2X1 NAND2X1_1904 ( .A(wSelec[2]), .B(_202_), .Y(_203_) );
	NOR2X1 NOR2X1_1078 ( .A(_203_), .B(_196_), .Y(_204_) );
	NAND2X1 NAND2X1_1905 ( .A(wData[24]), .B(_204_), .Y(_205_) );
	INVX1 INVX1_1164 ( .A(wSelec[3]), .Y(_206_) );
	NAND2X1 NAND2X1_1906 ( .A(_206_), .B(_195_), .Y(_207_) );
	NOR2X1 NOR2X1_1079 ( .A(_194_), .B(_207_), .Y(_208_) );
	NAND2X1 NAND2X1_1907 ( .A(wSelec[2]), .B(wSelec[1]), .Y(_209_) );
	NOR2X1 NOR2X1_1080 ( .A(_209_), .B(_196_), .Y(_210_) );
	AOI22X1 AOI22X1_1438 ( .A(_210_), .B(wData[28]), .C(wData[4]), .D(_208_), .Y(_211_) );
	NAND3X1 NAND3X1_509 ( .A(_205_), .B(_211_), .C(_201_), .Y(_212_) );
	NAND2X1 NAND2X1_1908 ( .A(wSelec[4]), .B(_206_), .Y(_213_) );
	NOR2X1 NOR2X1_1081 ( .A(_213_), .B(_199_), .Y(_214_) );
	NAND2X1 NAND2X1_1909 ( .A(wData[32]), .B(_214_), .Y(_215_) );
	NAND2X1 NAND2X1_1910 ( .A(wSelec[3]), .B(wSelec[4]), .Y(_216_) );
	NOR2X1 NOR2X1_1082 ( .A(_216_), .B(_203_), .Y(_217_) );
	NOR2X1 NOR2X1_1083 ( .A(_216_), .B(_194_), .Y(_218_) );
	AOI22X1 AOI22X1_1439 ( .A(_217_), .B(wData[56]), .C(wData[52]), .D(_218_), .Y(_219_) );
	NOR2X1 NOR2X1_1084 ( .A(_209_), .B(_216_), .Y(_220_) );
	NOR2X1 NOR2X1_1085 ( .A(_209_), .B(_213_), .Y(_221_) );
	AOI22X1 AOI22X1_1440 ( .A(wData[60]), .B(_220_), .C(_221_), .D(wData[44]), .Y(_222_) );
	NAND3X1 NAND3X1_510 ( .A(_215_), .B(_222_), .C(_219_), .Y(_223_) );
	NOR2X1 NOR2X1_1086 ( .A(_203_), .B(_213_), .Y(_224_) );
	NAND2X1 NAND2X1_1911 ( .A(wData[40]), .B(_224_), .Y(_225_) );
	NOR2X1 NOR2X1_1087 ( .A(_213_), .B(_194_), .Y(_226_) );
	NAND2X1 NAND2X1_1912 ( .A(wData[36]), .B(_226_), .Y(_227_) );
	NOR2X1 NOR2X1_1088 ( .A(_207_), .B(_199_), .Y(_228_) );
	NAND2X1 NAND2X1_1913 ( .A(wData[0]), .B(_228_), .Y(_229_) );
	NAND3X1 NAND3X1_511 ( .A(_225_), .B(_227_), .C(_229_), .Y(_230_) );
	INVX1 INVX1_1165 ( .A(wData[48]), .Y(_231_) );
	NOR2X1 NOR2X1_1089 ( .A(_206_), .B(_195_), .Y(_232_) );
	NAND2X1 NAND2X1_1914 ( .A(_198_), .B(_232_), .Y(_233_) );
	NOR2X1 NOR2X1_1090 ( .A(_203_), .B(_207_), .Y(_234_) );
	NOR2X1 NOR2X1_1091 ( .A(_209_), .B(_207_), .Y(_235_) );
	AOI22X1 AOI22X1_1441 ( .A(_234_), .B(wData[8]), .C(wData[12]), .D(_235_), .Y(_236_) );
	OAI21X1 OAI21X1_322 ( .A(_231_), .B(_233_), .C(_236_), .Y(_237_) );
	OR2X2 OR2X2_105 ( .A(_237_), .B(_230_), .Y(_238_) );
	NOR3X1 NOR3X1_787 ( .A(_212_), .B(_223_), .C(_238_), .Y(_239_) );
	AND2X2 AND2X2_200 ( .A(_239_), .B(_3_), .Y(_240_) );
	AOI21X1 AOI21X1_217 ( .A(_94_), .B(_192_), .C(_240_), .Y(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_0_) );
	INVX1 INVX1_1166 ( .A(_111_), .Y(_241_) );
	AOI21X1 AOI21X1_218 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_241_), .C(_3_), .Y(_242_) );
	AOI22X1 AOI22X1_1442 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_11_), .C(_27_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_243_) );
	AOI22X1 AOI22X1_1443 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_31_), .C(_37_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_244_) );
	NAND3X1 NAND3X1_512 ( .A(_242_), .B(_243_), .C(_244_), .Y(_245_) );
	INVX1 INVX1_1167 ( .A(_71_), .Y(_246_) );
	AOI22X1 AOI22X1_1444 ( .A(_96_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_246_), .Y(_247_) );
	AOI22X1 AOI22X1_1445 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_170_), .C(_49_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_248_) );
	INVX1 INVX1_1168 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_249_) );
	INVX1 INVX1_1169 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_250_) );
	OAI22X1 OAI22X1_247 ( .A(_249_), .B(_58_), .C(_56_), .D(_250_), .Y(_251_) );
	INVX1 INVX1_1170 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_252_) );
	NAND2X1 NAND2X1_1915 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_159_), .Y(_253_) );
	OAI21X1 OAI21X1_323 ( .A(_252_), .B(_64_), .C(_253_), .Y(_254_) );
	NOR2X1 NOR2X1_1092 ( .A(_251_), .B(_254_), .Y(_255_) );
	NAND3X1 NAND3X1_513 ( .A(_247_), .B(_248_), .C(_255_), .Y(_256_) );
	INVX1 INVX1_1171 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_257_) );
	NAND2X1 NAND2X1_1916 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_43_), .Y(_258_) );
	OAI21X1 OAI21X1_324 ( .A(_257_), .B(_73_), .C(_258_), .Y(_259_) );
	INVX1 INVX1_1172 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_260_) );
	INVX1 INVX1_1173 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_261_) );
	OAI22X1 OAI22X1_248 ( .A(_260_), .B(_79_), .C(_77_), .D(_261_), .Y(_262_) );
	NOR2X1 NOR2X1_1093 ( .A(_262_), .B(_259_), .Y(_263_) );
	AOI22X1 AOI22X1_1446 ( .A(_163_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_136_), .Y(_264_) );
	AND2X2 AND2X2_201 ( .A(_10_), .B(_25_), .Y(_265_) );
	AOI22X1 AOI22X1_1447 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_135_), .C(_265_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_266_) );
	NAND3X1 NAND3X1_514 ( .A(_264_), .B(_266_), .C(_263_), .Y(_267_) );
	NOR3X1 NOR3X1_788 ( .A(_267_), .B(_245_), .C(_256_), .Y(_268_) );
	INVX1 INVX1_1174 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_269_) );
	NAND2X1 NAND2X1_1917 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_98_), .Y(_270_) );
	OAI21X1 OAI21X1_325 ( .A(_100_), .B(_269_), .C(_270_), .Y(_271_) );
	AOI21X1 AOI21X1_219 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_147_), .C(_271_), .Y(_272_) );
	INVX1 INVX1_1175 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_273_) );
	INVX1 INVX1_1176 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_274_) );
	OAI22X1 OAI22X1_249 ( .A(_274_), .B(_106_), .C(_107_), .D(_273_), .Y(_275_) );
	INVX1 INVX1_1177 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_276_) );
	NAND2X1 NAND2X1_1918 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_116_), .Y(_277_) );
	OAI21X1 OAI21X1_326 ( .A(_17_), .B(_276_), .C(_277_), .Y(_278_) );
	NOR2X1 NOR2X1_1094 ( .A(_278_), .B(_275_), .Y(_279_) );
	INVX1 INVX1_1178 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_280_) );
	INVX1 INVX1_1179 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_281_) );
	OAI22X1 OAI22X1_250 ( .A(_112_), .B(_281_), .C(_118_), .D(_280_), .Y(_282_) );
	INVX1 INVX1_1180 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_283_) );
	NOR2X1 NOR2X1_1095 ( .A(_283_), .B(_123_), .Y(_284_) );
	INVX1 INVX1_1181 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_285_) );
	NOR2X1 NOR2X1_1096 ( .A(_285_), .B(_124_), .Y(_286_) );
	NOR3X1 NOR3X1_789 ( .A(_284_), .B(_282_), .C(_286_), .Y(_287_) );
	NAND3X1 NAND3X1_515 ( .A(_279_), .B(_272_), .C(_287_), .Y(_288_) );
	AOI22X1 AOI22X1_1448 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_128_), .C(_129_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_289_) );
	AOI22X1 AOI22X1_1449 ( .A(_131_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_132_), .Y(_290_) );
	NAND2X1 NAND2X1_1919 ( .A(_289_), .B(_290_), .Y(_291_) );
	AOI22X1 AOI22X1_1450 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_139_), .C(_138_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_292_) );
	AOI22X1 AOI22X1_1451 ( .A(_82_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_89_), .Y(_293_) );
	NAND2X1 NAND2X1_1920 ( .A(_292_), .B(_293_), .Y(_294_) );
	NOR2X1 NOR2X1_1097 ( .A(_291_), .B(_294_), .Y(_295_) );
	AOI22X1 AOI22X1_1452 ( .A(_143_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_144_), .Y(_296_) );
	AOI22X1 AOI22X1_1453 ( .A(_45_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_146_), .Y(_297_) );
	NAND2X1 NAND2X1_1921 ( .A(_296_), .B(_297_), .Y(_298_) );
	AOI22X1 AOI22X1_1454 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_150_), .C(_151_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_299_) );
	AOI22X1 AOI22X1_1455 ( .A(_153_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_154_), .Y(_300_) );
	NAND2X1 NAND2X1_1922 ( .A(_300_), .B(_299_), .Y(_301_) );
	NOR2X1 NOR2X1_1098 ( .A(_298_), .B(_301_), .Y(_302_) );
	NAND2X1 NAND2X1_1923 ( .A(_302_), .B(_295_), .Y(_303_) );
	AOI22X1 AOI22X1_1456 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_160_), .C(_61_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_304_) );
	AOI22X1 AOI22X1_1457 ( .A(_84_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_162_), .Y(_305_) );
	NAND2X1 NAND2X1_1924 ( .A(_304_), .B(_305_), .Y(_306_) );
	AOI22X1 AOI22X1_1458 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_51_), .C(_171_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_307_) );
	NAND2X1 NAND2X1_1925 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_166_), .Y(_308_) );
	NAND2X1 NAND2X1_1926 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_168_), .Y(_309_) );
	NAND3X1 NAND3X1_516 ( .A(_308_), .B(_309_), .C(_307_), .Y(_310_) );
	NOR2X1 NOR2X1_1099 ( .A(_310_), .B(_306_), .Y(_311_) );
	AOI22X1 AOI22X1_1459 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_175_), .C(_176_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_312_) );
	NAND2X1 NAND2X1_1927 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_178_), .Y(_313_) );
	NAND2X1 NAND2X1_1928 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_180_), .Y(_314_) );
	NAND3X1 NAND3X1_517 ( .A(_313_), .B(_314_), .C(_312_), .Y(_315_) );
	AOI22X1 AOI22X1_1460 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_184_), .C(_183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_316_) );
	AOI22X1 AOI22X1_1461 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_187_), .C(_186_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_317_) );
	NAND2X1 NAND2X1_1929 ( .A(_316_), .B(_317_), .Y(_318_) );
	NOR2X1 NOR2X1_1100 ( .A(_318_), .B(_315_), .Y(_319_) );
	NAND2X1 NAND2X1_1930 ( .A(_311_), .B(_319_), .Y(_320_) );
	NOR3X1 NOR3X1_790 ( .A(_303_), .B(_288_), .C(_320_), .Y(_321_) );
	AOI21X1 AOI21X1_220 ( .A(wData[21]), .B(_197_), .C(_2_), .Y(_322_) );
	AOI22X1 AOI22X1_1462 ( .A(_200_), .B(wData[17]), .C(wData[1]), .D(_228_), .Y(_323_) );
	AOI22X1 AOI22X1_1463 ( .A(_221_), .B(wData[45]), .C(wData[25]), .D(_204_), .Y(_324_) );
	NAND3X1 NAND3X1_518 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
	NAND3X1 NAND3X1_519 ( .A(wData[49]), .B(_198_), .C(_232_), .Y(_326_) );
	AOI22X1 AOI22X1_1464 ( .A(wData[61]), .B(_220_), .C(_208_), .D(wData[5]), .Y(_327_) );
	AND2X2 AND2X2_202 ( .A(_327_), .B(_326_), .Y(_328_) );
	AOI22X1 AOI22X1_1465 ( .A(_217_), .B(wData[57]), .C(wData[41]), .D(_224_), .Y(_329_) );
	AOI22X1 AOI22X1_1466 ( .A(wData[53]), .B(_218_), .C(_214_), .D(wData[33]), .Y(_330_) );
	AND2X2 AND2X2_203 ( .A(_330_), .B(_329_), .Y(_331_) );
	AOI22X1 AOI22X1_1467 ( .A(_234_), .B(wData[9]), .C(wData[13]), .D(_235_), .Y(_332_) );
	AOI22X1 AOI22X1_1468 ( .A(_210_), .B(wData[29]), .C(wData[37]), .D(_226_), .Y(_333_) );
	AND2X2 AND2X2_204 ( .A(_332_), .B(_333_), .Y(_334_) );
	NAND3X1 NAND3X1_520 ( .A(_328_), .B(_334_), .C(_331_), .Y(_335_) );
	NOR2X1 NOR2X1_1101 ( .A(_325_), .B(_335_), .Y(_336_) );
	AOI21X1 AOI21X1_221 ( .A(_268_), .B(_321_), .C(_336_), .Y(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_1_) );
	AOI21X1 AOI21X1_222 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_241_), .C(_3_), .Y(_337_) );
	INVX1 INVX1_1182 ( .A(_100_), .Y(_338_) );
	AOI22X1 AOI22X1_1469 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_11_), .C(_338_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_339_) );
	INVX1 INVX1_1183 ( .A(_112_), .Y(_340_) );
	AOI22X1 AOI22X1_1470 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_147_), .C(_340_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_341_) );
	NAND3X1 NAND3X1_521 ( .A(_341_), .B(_337_), .C(_339_), .Y(_342_) );
	AOI22X1 AOI22X1_1471 ( .A(_96_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_246_), .Y(_343_) );
	AOI22X1 AOI22X1_1472 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_45_), .C(_18_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_344_) );
	INVX1 INVX1_1184 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_345_) );
	NAND2X1 NAND2X1_1931 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_135_), .Y(_346_) );
	OAI21X1 OAI21X1_327 ( .A(_345_), .B(_107_), .C(_346_), .Y(_347_) );
	INVX1 INVX1_1185 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_348_) );
	NAND2X1 NAND2X1_1932 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_61_), .Y(_349_) );
	OAI21X1 OAI21X1_328 ( .A(_348_), .B(_64_), .C(_349_), .Y(_350_) );
	NOR2X1 NOR2X1_1102 ( .A(_347_), .B(_350_), .Y(_351_) );
	NAND3X1 NAND3X1_522 ( .A(_343_), .B(_344_), .C(_351_), .Y(_352_) );
	INVX1 INVX1_1186 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_353_) );
	NAND2X1 NAND2X1_1933 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_43_), .Y(_354_) );
	OAI21X1 OAI21X1_329 ( .A(_353_), .B(_73_), .C(_354_), .Y(_355_) );
	INVX1 INVX1_1187 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_356_) );
	INVX1 INVX1_1188 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_357_) );
	OAI22X1 OAI22X1_251 ( .A(_356_), .B(_79_), .C(_77_), .D(_357_), .Y(_358_) );
	NOR2X1 NOR2X1_1103 ( .A(_358_), .B(_355_), .Y(_359_) );
	AOI22X1 AOI22X1_1473 ( .A(_163_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_136_), .Y(_360_) );
	AND2X2 AND2X2_205 ( .A(_35_), .B(_57_), .Y(_361_) );
	AOI22X1 AOI22X1_1474 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_361_), .C(_265_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_362_) );
	NAND3X1 NAND3X1_523 ( .A(_360_), .B(_362_), .C(_359_), .Y(_363_) );
	NOR3X1 NOR3X1_791 ( .A(_363_), .B(_342_), .C(_352_), .Y(_364_) );
	INVX1 INVX1_1189 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_365_) );
	NOR3X1 NOR3X1_792 ( .A(_365_), .B(_30_), .C(_29_), .Y(_366_) );
	AND2X2 AND2X2_206 ( .A(_51_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_367_) );
	AND2X2 AND2X2_207 ( .A(_171_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_368_) );
	NOR3X1 NOR3X1_793 ( .A(_368_), .B(_367_), .C(_366_), .Y(_369_) );
	INVX1 INVX1_1190 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_370_) );
	INVX1 INVX1_1191 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_371_) );
	OAI22X1 OAI22X1_252 ( .A(_371_), .B(_106_), .C(_56_), .D(_370_), .Y(_372_) );
	INVX1 INVX1_1192 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_373_) );
	INVX1 INVX1_1193 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_374_) );
	NAND2X1 NAND2X1_1934 ( .A(_47_), .B(_48_), .Y(_375_) );
	OAI22X1 OAI22X1_253 ( .A(_375_), .B(_374_), .C(_373_), .D(_26_), .Y(_376_) );
	NOR2X1 NOR2X1_1104 ( .A(_372_), .B(_376_), .Y(_377_) );
	INVX1 INVX1_1194 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_378_) );
	NOR3X1 NOR3X1_794 ( .A(_7_), .B(_24_), .C(_15_), .Y(_379_) );
	NAND2X1 NAND2X1_1935 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_379_), .Y(_380_) );
	OAI21X1 OAI21X1_330 ( .A(_36_), .B(_378_), .C(_380_), .Y(_381_) );
	INVX1 INVX1_1195 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_382_) );
	INVX1 INVX1_1196 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_383_) );
	OAI22X1 OAI22X1_254 ( .A(_123_), .B(_383_), .C(_382_), .D(_124_), .Y(_384_) );
	NOR2X1 NOR2X1_1105 ( .A(_381_), .B(_384_), .Y(_385_) );
	NAND3X1 NAND3X1_524 ( .A(_369_), .B(_385_), .C(_377_), .Y(_386_) );
	AOI22X1 AOI22X1_1475 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_128_), .C(_129_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_387_) );
	AOI22X1 AOI22X1_1476 ( .A(_131_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_132_), .Y(_388_) );
	NAND2X1 NAND2X1_1936 ( .A(_387_), .B(_388_), .Y(_389_) );
	AOI22X1 AOI22X1_1477 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_139_), .C(_138_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_390_) );
	AOI22X1 AOI22X1_1478 ( .A(_82_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_89_), .Y(_391_) );
	NAND2X1 NAND2X1_1937 ( .A(_390_), .B(_391_), .Y(_392_) );
	NOR2X1 NOR2X1_1106 ( .A(_389_), .B(_392_), .Y(_393_) );
	AOI22X1 AOI22X1_1479 ( .A(_143_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_144_), .Y(_394_) );
	AOI22X1 AOI22X1_1480 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_170_), .C(_146_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_395_) );
	NAND2X1 NAND2X1_1938 ( .A(_395_), .B(_394_), .Y(_396_) );
	AOI22X1 AOI22X1_1481 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_150_), .C(_151_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_397_) );
	AOI22X1 AOI22X1_1482 ( .A(_153_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_154_), .Y(_398_) );
	NAND2X1 NAND2X1_1939 ( .A(_398_), .B(_397_), .Y(_399_) );
	NOR2X1 NOR2X1_1107 ( .A(_396_), .B(_399_), .Y(_400_) );
	NAND2X1 NAND2X1_1940 ( .A(_400_), .B(_393_), .Y(_401_) );
	AOI22X1 AOI22X1_1483 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_160_), .C(_159_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_402_) );
	AOI22X1 AOI22X1_1484 ( .A(_84_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_162_), .Y(_403_) );
	NAND2X1 NAND2X1_1941 ( .A(_402_), .B(_403_), .Y(_404_) );
	AOI22X1 AOI22X1_1485 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_168_), .C(_166_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_405_) );
	AOI22X1 AOI22X1_1486 ( .A(_98_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_116_), .Y(_406_) );
	NAND2X1 NAND2X1_1942 ( .A(_406_), .B(_405_), .Y(_407_) );
	NOR2X1 NOR2X1_1108 ( .A(_407_), .B(_404_), .Y(_408_) );
	AOI22X1 AOI22X1_1487 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_175_), .C(_176_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_409_) );
	NAND2X1 NAND2X1_1943 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_178_), .Y(_410_) );
	NAND2X1 NAND2X1_1944 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_180_), .Y(_411_) );
	NAND3X1 NAND3X1_525 ( .A(_410_), .B(_411_), .C(_409_), .Y(_412_) );
	AOI22X1 AOI22X1_1488 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_184_), .C(_183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_413_) );
	AOI22X1 AOI22X1_1489 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_187_), .C(_186_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_414_) );
	NAND2X1 NAND2X1_1945 ( .A(_413_), .B(_414_), .Y(_415_) );
	NOR2X1 NOR2X1_1109 ( .A(_415_), .B(_412_), .Y(_416_) );
	NAND2X1 NAND2X1_1946 ( .A(_408_), .B(_416_), .Y(_417_) );
	NOR3X1 NOR3X1_795 ( .A(_401_), .B(_386_), .C(_417_), .Y(_418_) );
	AOI22X1 AOI22X1_1490 ( .A(_224_), .B(wData[42]), .C(wData[38]), .D(_226_), .Y(_419_) );
	AOI22X1 AOI22X1_1491 ( .A(_221_), .B(wData[46]), .C(_228_), .D(wData[2]), .Y(_420_) );
	NAND2X1 NAND2X1_1947 ( .A(_419_), .B(_420_), .Y(_421_) );
	AOI21X1 AOI21X1_223 ( .A(wData[34]), .B(_214_), .C(_421_), .Y(_422_) );
	INVX1 INVX1_1197 ( .A(wData[50]), .Y(_423_) );
	AOI22X1 AOI22X1_1492 ( .A(_234_), .B(wData[10]), .C(wData[14]), .D(_235_), .Y(_424_) );
	OAI21X1 OAI21X1_331 ( .A(_423_), .B(_233_), .C(_424_), .Y(_425_) );
	AOI22X1 AOI22X1_1493 ( .A(_197_), .B(wData[22]), .C(wData[18]), .D(_200_), .Y(_426_) );
	NAND2X1 NAND2X1_1948 ( .A(wData[26]), .B(_204_), .Y(_427_) );
	AOI22X1 AOI22X1_1494 ( .A(_210_), .B(wData[30]), .C(wData[6]), .D(_208_), .Y(_428_) );
	NAND3X1 NAND3X1_526 ( .A(_427_), .B(_428_), .C(_426_), .Y(_429_) );
	NOR2X1 NOR2X1_1110 ( .A(_425_), .B(_429_), .Y(_430_) );
	NAND2X1 NAND2X1_1949 ( .A(wData[58]), .B(_217_), .Y(_431_) );
	NAND2X1 NAND2X1_1950 ( .A(wData[54]), .B(_218_), .Y(_432_) );
	NAND2X1 NAND2X1_1951 ( .A(_431_), .B(_432_), .Y(_433_) );
	AOI21X1 AOI21X1_224 ( .A(wData[62]), .B(_220_), .C(_433_), .Y(_434_) );
	NAND3X1 NAND3X1_527 ( .A(_422_), .B(_434_), .C(_430_), .Y(_435_) );
	NOR2X1 NOR2X1_1111 ( .A(_2_), .B(_435_), .Y(_436_) );
	AOI21X1 AOI21X1_225 ( .A(_364_), .B(_418_), .C(_436_), .Y(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_2_) );
	AOI21X1 AOI21X1_226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_246_), .C(_3_), .Y(_437_) );
	AOI22X1 AOI22X1_1495 ( .A(_18_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_338_), .Y(_438_) );
	AOI22X1 AOI22X1_1496 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_340_), .C(_96_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_439_) );
	NAND3X1 NAND3X1_528 ( .A(_439_), .B(_437_), .C(_438_), .Y(_440_) );
	AOI22X1 AOI22X1_1497 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_45_), .C(_43_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_441_) );
	AOI22X1 AOI22X1_1498 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_116_), .C(_241_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_442_) );
	INVX1 INVX1_1198 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_443_) );
	INVX1 INVX1_1199 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_444_) );
	OAI22X1 OAI22X1_255 ( .A(_443_), .B(_58_), .C(_107_), .D(_444_), .Y(_445_) );
	INVX1 INVX1_1200 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_446_) );
	NAND2X1 NAND2X1_1952 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_159_), .Y(_447_) );
	OAI21X1 OAI21X1_332 ( .A(_446_), .B(_64_), .C(_447_), .Y(_448_) );
	NOR2X1 NOR2X1_1112 ( .A(_445_), .B(_448_), .Y(_449_) );
	NAND3X1 NAND3X1_529 ( .A(_441_), .B(_442_), .C(_449_), .Y(_450_) );
	AND2X2 AND2X2_208 ( .A(_72_), .B(_6_), .Y(_451_) );
	AOI22X1 AOI22X1_1499 ( .A(_11_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_451_), .Y(_452_) );
	AND2X2 AND2X2_209 ( .A(_70_), .B(_35_), .Y(_453_) );
	AND2X2 AND2X2_210 ( .A(_78_), .B(_35_), .Y(_454_) );
	AOI22X1 AOI22X1_1500 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_454_), .C(_453_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_455_) );
	NAND2X1 NAND2X1_1953 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__3_), .B(_163_), .Y(_456_) );
	NAND2X1 NAND2X1_1954 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__3_), .B(_136_), .Y(_457_) );
	NAND2X1 NAND2X1_1955 ( .A(_456_), .B(_457_), .Y(_458_) );
	INVX1 INVX1_1201 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__3_), .Y(_459_) );
	NAND2X1 NAND2X1_1956 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__3_), .B(_135_), .Y(_460_) );
	OAI21X1 OAI21X1_333 ( .A(_459_), .B(_88_), .C(_460_), .Y(_461_) );
	NOR2X1 NOR2X1_1113 ( .A(_458_), .B(_461_), .Y(_462_) );
	NAND3X1 NAND3X1_530 ( .A(_452_), .B(_455_), .C(_462_), .Y(_463_) );
	NOR3X1 NOR3X1_796 ( .A(_450_), .B(_440_), .C(_463_), .Y(_464_) );
	INVX1 INVX1_1202 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__3_), .Y(_465_) );
	NAND2X1 NAND2X1_1957 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__3_), .B(_51_), .Y(_466_) );
	OAI21X1 OAI21X1_334 ( .A(_56_), .B(_465_), .C(_466_), .Y(_467_) );
	AOI21X1 AOI21X1_227 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__3_), .B(_31_), .C(_467_), .Y(_468_) );
	INVX1 INVX1_1203 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__3_), .Y(_469_) );
	INVX1 INVX1_1204 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__3_), .Y(_470_) );
	OAI22X1 OAI22X1_256 ( .A(_375_), .B(_470_), .C(_469_), .D(_26_), .Y(_471_) );
	INVX1 INVX1_1205 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__3_), .Y(_472_) );
	NAND2X1 NAND2X1_1958 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__3_), .B(_171_), .Y(_473_) );
	OAI21X1 OAI21X1_335 ( .A(_36_), .B(_472_), .C(_473_), .Y(_474_) );
	NOR2X1 NOR2X1_1114 ( .A(_474_), .B(_471_), .Y(_475_) );
	INVX1 INVX1_1206 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__3_), .Y(_476_) );
	INVX1 INVX1_1207 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__3_), .Y(_477_) );
	OAI22X1 OAI22X1_257 ( .A(_123_), .B(_477_), .C(_476_), .D(_124_), .Y(_478_) );
	INVX1 INVX1_1208 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__3_), .Y(_479_) );
	NAND2X1 NAND2X1_1959 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__3_), .B(_170_), .Y(_480_) );
	OAI21X1 OAI21X1_336 ( .A(_479_), .B(_106_), .C(_480_), .Y(_481_) );
	NOR2X1 NOR2X1_1115 ( .A(_481_), .B(_478_), .Y(_482_) );
	NAND3X1 NAND3X1_531 ( .A(_468_), .B(_482_), .C(_475_), .Y(_483_) );
	AOI22X1 AOI22X1_1501 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__3_), .B(_128_), .C(_129_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__3_), .Y(_484_) );
	AOI22X1 AOI22X1_1502 ( .A(_131_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__3_), .D(_132_), .Y(_485_) );
	NAND2X1 NAND2X1_1960 ( .A(_484_), .B(_485_), .Y(_486_) );
	AOI22X1 AOI22X1_1503 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__3_), .B(_139_), .C(_138_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__3_), .Y(_487_) );
	AOI22X1 AOI22X1_1504 ( .A(_82_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__3_), .D(_89_), .Y(_488_) );
	NAND2X1 NAND2X1_1961 ( .A(_487_), .B(_488_), .Y(_489_) );
	NOR2X1 NOR2X1_1116 ( .A(_486_), .B(_489_), .Y(_490_) );
	AOI22X1 AOI22X1_1505 ( .A(_143_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__3_), .D(_144_), .Y(_491_) );
	AOI22X1 AOI22X1_1506 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__3_), .B(_379_), .C(_146_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__3_), .Y(_492_) );
	NAND2X1 NAND2X1_1962 ( .A(_492_), .B(_491_), .Y(_493_) );
	AOI22X1 AOI22X1_1507 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__3_), .B(_150_), .C(_151_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__3_), .Y(_494_) );
	AOI22X1 AOI22X1_1508 ( .A(_153_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__3_), .D(_154_), .Y(_495_) );
	NAND2X1 NAND2X1_1963 ( .A(_495_), .B(_494_), .Y(_496_) );
	NOR2X1 NOR2X1_1117 ( .A(_493_), .B(_496_), .Y(_497_) );
	NAND2X1 NAND2X1_1964 ( .A(_497_), .B(_490_), .Y(_498_) );
	AOI22X1 AOI22X1_1509 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__3_), .B(_160_), .C(_61_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__3_), .Y(_499_) );
	AOI22X1 AOI22X1_1510 ( .A(_84_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__3_), .D(_162_), .Y(_500_) );
	NAND2X1 NAND2X1_1965 ( .A(_499_), .B(_500_), .Y(_501_) );
	AOI22X1 AOI22X1_1511 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__3_), .B(_168_), .C(_166_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__3_), .Y(_502_) );
	AOI22X1 AOI22X1_1512 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__3_), .B(_98_), .C(_147_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__3_), .Y(_503_) );
	NAND2X1 NAND2X1_1966 ( .A(_503_), .B(_502_), .Y(_504_) );
	NOR2X1 NOR2X1_1118 ( .A(_504_), .B(_501_), .Y(_505_) );
	AOI22X1 AOI22X1_1513 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__3_), .B(_175_), .C(_176_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__3_), .Y(_506_) );
	NAND2X1 NAND2X1_1967 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__3_), .B(_178_), .Y(_507_) );
	NAND2X1 NAND2X1_1968 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__3_), .B(_180_), .Y(_508_) );
	NAND3X1 NAND3X1_532 ( .A(_507_), .B(_508_), .C(_506_), .Y(_509_) );
	AOI22X1 AOI22X1_1514 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__3_), .B(_184_), .C(_183_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__3_), .Y(_510_) );
	AOI22X1 AOI22X1_1515 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__3_), .B(_187_), .C(_186_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__3_), .Y(_511_) );
	NAND2X1 NAND2X1_1969 ( .A(_510_), .B(_511_), .Y(_512_) );
	NOR2X1 NOR2X1_1119 ( .A(_512_), .B(_509_), .Y(_513_) );
	NAND2X1 NAND2X1_1970 ( .A(_505_), .B(_513_), .Y(_514_) );
	NOR3X1 NOR3X1_797 ( .A(_498_), .B(_483_), .C(_514_), .Y(_515_) );
	NAND2X1 NAND2X1_1971 ( .A(wData[59]), .B(_217_), .Y(_516_) );
	OAI21X1 OAI21X1_337 ( .A(_1_), .B(wBusy_bF_buf4), .C(_516_), .Y(_517_) );
	NAND2X1 NAND2X1_1972 ( .A(wData[7]), .B(_208_), .Y(_518_) );
	NAND2X1 NAND2X1_1973 ( .A(wData[55]), .B(_218_), .Y(_519_) );
	AOI22X1 AOI22X1_1516 ( .A(wData[63]), .B(_220_), .C(_210_), .D(wData[31]), .Y(_520_) );
	NAND3X1 NAND3X1_533 ( .A(_518_), .B(_519_), .C(_520_), .Y(_521_) );
	OR2X2 OR2X2_106 ( .A(_521_), .B(_517_), .Y(_522_) );
	INVX1 INVX1_1209 ( .A(wData[51]), .Y(_523_) );
	NAND2X1 NAND2X1_1974 ( .A(wData[47]), .B(_221_), .Y(_524_) );
	OAI21X1 OAI21X1_338 ( .A(_523_), .B(_233_), .C(_524_), .Y(_525_) );
	AOI21X1 AOI21X1_228 ( .A(wData[3]), .B(_228_), .C(_525_), .Y(_526_) );
	AOI22X1 AOI22X1_1517 ( .A(_234_), .B(wData[11]), .C(wData[15]), .D(_235_), .Y(_527_) );
	AOI22X1 AOI22X1_1518 ( .A(_197_), .B(wData[23]), .C(wData[27]), .D(_204_), .Y(_528_) );
	AND2X2 AND2X2_211 ( .A(_527_), .B(_528_), .Y(_529_) );
	NAND2X1 NAND2X1_1975 ( .A(wData[39]), .B(_226_), .Y(_530_) );
	NAND2X1 NAND2X1_1976 ( .A(wData[43]), .B(_224_), .Y(_531_) );
	NAND2X1 NAND2X1_1977 ( .A(_530_), .B(_531_), .Y(_532_) );
	NAND2X1 NAND2X1_1978 ( .A(wData[19]), .B(_200_), .Y(_533_) );
	NAND2X1 NAND2X1_1979 ( .A(wData[35]), .B(_214_), .Y(_534_) );
	NAND2X1 NAND2X1_1980 ( .A(_533_), .B(_534_), .Y(_535_) );
	NOR2X1 NOR2X1_1120 ( .A(_532_), .B(_535_), .Y(_536_) );
	NAND3X1 NAND3X1_534 ( .A(_529_), .B(_526_), .C(_536_), .Y(_537_) );
	NOR2X1 NOR2X1_1121 ( .A(_522_), .B(_537_), .Y(_538_) );
	AOI21X1 AOI21X1_229 ( .A(_464_), .B(_515_), .C(_538_), .Y(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_r_3_) );
	INVX1 INVX1_1210 ( .A(wSelec[11]), .Y(_539_) );
	NOR2X1 NOR2X1_1122 ( .A(wBusy_bF_buf3), .B(_539_), .Y(_540_) );
	INVX1 INVX1_1211 ( .A(_540_), .Y(_541_) );
	INVX1 INVX1_1212 ( .A(wSelec[21]), .Y(_542_) );
	NAND2X1 NAND2X1_1981 ( .A(wSelec[20]), .B(_542_), .Y(_543_) );
	INVX2 INVX2_31 ( .A(_543_), .Y(_544_) );
	OR2X2 OR2X2_107 ( .A(wSelec[17]), .B(wSelec[16]), .Y(_545_) );
	INVX1 INVX1_1213 ( .A(wSelec[19]), .Y(_546_) );
	NAND2X1 NAND2X1_1982 ( .A(wSelec[18]), .B(_546_), .Y(_547_) );
	NOR2X1 NOR2X1_1123 ( .A(_545_), .B(_547_), .Y(_548_) );
	AND2X2 AND2X2_212 ( .A(_548_), .B(_544_), .Y(_549_) );
	AOI21X1 AOI21X1_230 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__0_), .B(_549_), .C(_541_), .Y(_550_) );
	INVX1 INVX1_1214 ( .A(wSelec[17]), .Y(_551_) );
	NAND2X1 NAND2X1_1983 ( .A(wSelec[16]), .B(_551_), .Y(_552_) );
	OR2X2 OR2X2_108 ( .A(wSelec[18]), .B(wSelec[19]), .Y(_553_) );
	NOR2X1 NOR2X1_1124 ( .A(_553_), .B(_552_), .Y(_554_) );
	NAND2X1 NAND2X1_1984 ( .A(_544_), .B(_554_), .Y(_555_) );
	INVX1 INVX1_1215 ( .A(_555_), .Y(_556_) );
	INVX1 INVX1_1216 ( .A(wSelec[16]), .Y(_557_) );
	NAND2X1 NAND2X1_1985 ( .A(wSelec[17]), .B(_557_), .Y(_558_) );
	INVX1 INVX1_1217 ( .A(wSelec[18]), .Y(_559_) );
	NAND2X1 NAND2X1_1986 ( .A(wSelec[19]), .B(_559_), .Y(_560_) );
	NOR2X1 NOR2X1_1125 ( .A(_558_), .B(_560_), .Y(_561_) );
	NAND2X1 NAND2X1_1987 ( .A(wSelec[20]), .B(wSelec[21]), .Y(_562_) );
	INVX1 INVX1_1218 ( .A(_562_), .Y(_563_) );
	NAND2X1 NAND2X1_1988 ( .A(_563_), .B(_561_), .Y(_564_) );
	INVX1 INVX1_1219 ( .A(_564_), .Y(_565_) );
	AOI22X1 AOI22X1_1519 ( .A(_556_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__0_), .D(_565_), .Y(_566_) );
	OR2X2 OR2X2_109 ( .A(_552_), .B(_553_), .Y(_567_) );
	OR2X2 OR2X2_110 ( .A(wSelec[20]), .B(wSelec[21]), .Y(_568_) );
	NOR2X1 NOR2X1_1126 ( .A(_568_), .B(_567_), .Y(_569_) );
	NOR2X1 NOR2X1_1127 ( .A(_547_), .B(_552_), .Y(_570_) );
	INVX1 INVX1_1220 ( .A(wSelec[20]), .Y(_571_) );
	NAND2X1 NAND2X1_1989 ( .A(wSelec[21]), .B(_571_), .Y(_572_) );
	INVX2 INVX2_32 ( .A(_572_), .Y(_573_) );
	NAND2X1 NAND2X1_1990 ( .A(_573_), .B(_570_), .Y(_574_) );
	INVX1 INVX1_1221 ( .A(_574_), .Y(_575_) );
	AOI22X1 AOI22X1_1520 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__0_), .B(_569_), .C(_575_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__0_), .Y(_576_) );
	NAND3X1 NAND3X1_535 ( .A(_550_), .B(_576_), .C(_566_), .Y(_577_) );
	NOR2X1 NOR2X1_1128 ( .A(wSelec[17]), .B(wSelec[16]), .Y(_578_) );
	NOR2X1 NOR2X1_1129 ( .A(wSelec[18]), .B(wSelec[19]), .Y(_579_) );
	NAND2X1 NAND2X1_1991 ( .A(_578_), .B(_579_), .Y(_580_) );
	NOR2X1 NOR2X1_1130 ( .A(_543_), .B(_580_), .Y(_581_) );
	NAND2X1 NAND2X1_1992 ( .A(wSelec[17]), .B(wSelec[16]), .Y(_582_) );
	NOR3X1 NOR3X1_798 ( .A(_553_), .B(_582_), .C(_543_), .Y(_583_) );
	AOI22X1 AOI22X1_1521 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__0_), .B(_583_), .C(_581_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__0_), .Y(_584_) );
	INVX1 INVX1_1222 ( .A(_568_), .Y(_585_) );
	NOR2X1 NOR2X1_1131 ( .A(_553_), .B(_558_), .Y(_586_) );
	AND2X2 AND2X2_213 ( .A(_586_), .B(_585_), .Y(_587_) );
	NAND2X1 NAND2X1_1993 ( .A(wSelec[18]), .B(wSelec[19]), .Y(_588_) );
	NOR3X1 NOR3X1_799 ( .A(_562_), .B(_582_), .C(_588_), .Y(_589_) );
	AOI22X1 AOI22X1_1522 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__0_), .B(_589_), .C(_587_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__0_), .Y(_590_) );
	INVX1 INVX1_1223 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__0_), .Y(_591_) );
	INVX1 INVX1_1224 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__0_), .Y(_592_) );
	NOR2X1 NOR2X1_1132 ( .A(_552_), .B(_560_), .Y(_593_) );
	NAND2X1 NAND2X1_1994 ( .A(_563_), .B(_593_), .Y(_594_) );
	NOR2X1 NOR2X1_1133 ( .A(_582_), .B(_588_), .Y(_595_) );
	NAND2X1 NAND2X1_1995 ( .A(_595_), .B(_573_), .Y(_596_) );
	OAI22X1 OAI22X1_258 ( .A(_591_), .B(_596_), .C(_594_), .D(_592_), .Y(_597_) );
	INVX1 INVX1_1225 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__0_), .Y(_598_) );
	NOR3X1 NOR3X1_800 ( .A(_543_), .B(_558_), .C(_560_), .Y(_599_) );
	NAND2X1 NAND2X1_1996 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__0_), .B(_599_), .Y(_600_) );
	NOR2X1 NOR2X1_1134 ( .A(_582_), .B(_547_), .Y(_601_) );
	NAND2X1 NAND2X1_1997 ( .A(_573_), .B(_601_), .Y(_602_) );
	OAI21X1 OAI21X1_339 ( .A(_598_), .B(_602_), .C(_600_), .Y(_603_) );
	NOR2X1 NOR2X1_1135 ( .A(_597_), .B(_603_), .Y(_604_) );
	NAND3X1 NAND3X1_536 ( .A(_584_), .B(_590_), .C(_604_), .Y(_605_) );
	INVX1 INVX1_1226 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__0_), .Y(_606_) );
	INVX1 INVX1_1227 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__0_), .Y(_607_) );
	NOR2X1 NOR2X1_1136 ( .A(_547_), .B(_558_), .Y(_608_) );
	NAND2X1 NAND2X1_1998 ( .A(_544_), .B(_608_), .Y(_609_) );
	NOR2X1 NOR2X1_1137 ( .A(_545_), .B(_560_), .Y(_610_) );
	NAND2X1 NAND2X1_1999 ( .A(_544_), .B(_610_), .Y(_611_) );
	OAI22X1 OAI22X1_259 ( .A(_611_), .B(_606_), .C(_607_), .D(_609_), .Y(_612_) );
	INVX1 INVX1_1228 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__0_), .Y(_613_) );
	INVX1 INVX1_1229 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__0_), .Y(_614_) );
	NAND2X1 NAND2X1_2000 ( .A(_573_), .B(_608_), .Y(_615_) );
	NOR2X1 NOR2X1_1138 ( .A(_582_), .B(_553_), .Y(_616_) );
	NAND2X1 NAND2X1_2001 ( .A(_573_), .B(_616_), .Y(_617_) );
	OAI22X1 OAI22X1_260 ( .A(_613_), .B(_617_), .C(_615_), .D(_614_), .Y(_618_) );
	NOR2X1 NOR2X1_1139 ( .A(_618_), .B(_612_), .Y(_619_) );
	NOR3X1 NOR3X1_801 ( .A(_552_), .B(_588_), .C(_572_), .Y(_620_) );
	NAND2X1 NAND2X1_2002 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__0_), .B(_620_), .Y(_621_) );
	NOR3X1 NOR3X1_802 ( .A(_560_), .B(_582_), .C(_572_), .Y(_622_) );
	NAND2X1 NAND2X1_2003 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__0_), .B(_622_), .Y(_623_) );
	NAND2X1 NAND2X1_2004 ( .A(_621_), .B(_623_), .Y(_624_) );
	INVX1 INVX1_1230 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__0_), .Y(_625_) );
	NAND2X1 NAND2X1_2005 ( .A(_563_), .B(_548_), .Y(_626_) );
	NOR3X1 NOR3X1_803 ( .A(_558_), .B(_560_), .C(_572_), .Y(_627_) );
	NAND2X1 NAND2X1_2006 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__0_), .B(_627_), .Y(_628_) );
	OAI21X1 OAI21X1_340 ( .A(_625_), .B(_626_), .C(_628_), .Y(_629_) );
	NOR2X1 NOR2X1_1140 ( .A(_624_), .B(_629_), .Y(_630_) );
	NAND2X1 NAND2X1_2007 ( .A(_619_), .B(_630_), .Y(_631_) );
	NOR3X1 NOR3X1_804 ( .A(_577_), .B(_631_), .C(_605_), .Y(_632_) );
	NAND2X1 NAND2X1_2008 ( .A(_544_), .B(_601_), .Y(_633_) );
	INVX1 INVX1_1231 ( .A(_633_), .Y(_634_) );
	INVX1 INVX1_1232 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__0_), .Y(_635_) );
	NOR3X1 NOR3X1_805 ( .A(_545_), .B(_568_), .C(_547_), .Y(_636_) );
	NAND2X1 NAND2X1_2009 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__0_), .B(_636_), .Y(_637_) );
	NAND2X1 NAND2X1_2010 ( .A(_585_), .B(_608_), .Y(_638_) );
	OAI21X1 OAI21X1_341 ( .A(_638_), .B(_635_), .C(_637_), .Y(_639_) );
	AOI21X1 AOI21X1_231 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__0_), .B(_634_), .C(_639_), .Y(_640_) );
	INVX1 INVX1_1233 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__0_), .Y(_641_) );
	INVX1 INVX1_1234 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__0_), .Y(_642_) );
	NOR2X1 NOR2X1_1141 ( .A(_588_), .B(_545_), .Y(_643_) );
	NAND2X1 NAND2X1_2011 ( .A(_544_), .B(_643_), .Y(_644_) );
	NAND2X1 NAND2X1_2012 ( .A(_585_), .B(_570_), .Y(_645_) );
	OAI22X1 OAI22X1_261 ( .A(_642_), .B(_644_), .C(_645_), .D(_641_), .Y(_646_) );
	INVX1 INVX1_1235 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__0_), .Y(_647_) );
	INVX1 INVX1_1236 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__0_), .Y(_648_) );
	NAND2X1 NAND2X1_2013 ( .A(_544_), .B(_570_), .Y(_649_) );
	NAND2X1 NAND2X1_2014 ( .A(_585_), .B(_616_), .Y(_650_) );
	OAI22X1 OAI22X1_262 ( .A(_647_), .B(_650_), .C(_649_), .D(_648_), .Y(_651_) );
	NOR2X1 NOR2X1_1142 ( .A(_646_), .B(_651_), .Y(_652_) );
	INVX1 INVX1_1237 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__0_), .Y(_653_) );
	NOR3X1 NOR3X1_806 ( .A(_568_), .B(_582_), .C(_547_), .Y(_654_) );
	NAND2X1 NAND2X1_2015 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__0_), .B(_654_), .Y(_655_) );
	OR2X2 OR2X2_111 ( .A(_580_), .B(_562_), .Y(_656_) );
	OAI21X1 OAI21X1_342 ( .A(_653_), .B(_656_), .C(_655_), .Y(_657_) );
	INVX1 INVX1_1238 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__0_), .Y(_658_) );
	INVX1 INVX1_1239 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__0_), .Y(_659_) );
	NOR2X1 NOR2X1_1143 ( .A(_588_), .B(_558_), .Y(_660_) );
	NAND2X1 NAND2X1_2016 ( .A(_544_), .B(_660_), .Y(_661_) );
	NAND2X1 NAND2X1_2017 ( .A(_563_), .B(_554_), .Y(_662_) );
	OAI22X1 OAI22X1_263 ( .A(_661_), .B(_659_), .C(_658_), .D(_662_), .Y(_663_) );
	NOR2X1 NOR2X1_1144 ( .A(_657_), .B(_663_), .Y(_664_) );
	NAND3X1 NAND3X1_537 ( .A(_640_), .B(_664_), .C(_652_), .Y(_665_) );
	NOR3X1 NOR3X1_807 ( .A(_545_), .B(_553_), .C(_568_), .Y(_666_) );
	NOR3X1 NOR3X1_808 ( .A(_562_), .B(_588_), .C(_552_), .Y(_667_) );
	AOI22X1 AOI22X1_1523 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__0_), .B(_666_), .C(_667_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__0_), .Y(_668_) );
	NOR3X1 NOR3X1_809 ( .A(_562_), .B(_588_), .C(_558_), .Y(_669_) );
	NOR3X1 NOR3X1_810 ( .A(_562_), .B(_582_), .C(_560_), .Y(_670_) );
	AOI22X1 AOI22X1_1524 ( .A(_669_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__0_), .D(_670_), .Y(_671_) );
	NAND2X1 NAND2X1_2018 ( .A(_668_), .B(_671_), .Y(_672_) );
	NOR3X1 NOR3X1_811 ( .A(_560_), .B(_545_), .C(_572_), .Y(_673_) );
	NOR3X1 NOR3X1_812 ( .A(_552_), .B(_560_), .C(_572_), .Y(_674_) );
	AOI22X1 AOI22X1_1525 ( .A(_673_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__0_), .D(_674_), .Y(_675_) );
	NOR3X1 NOR3X1_813 ( .A(_543_), .B(_588_), .C(_552_), .Y(_676_) );
	NOR3X1 NOR3X1_814 ( .A(_582_), .B(_588_), .C(_543_), .Y(_677_) );
	AOI22X1 AOI22X1_1526 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__0_), .B(_677_), .C(_676_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__0_), .Y(_678_) );
	NAND2X1 NAND2X1_2019 ( .A(_678_), .B(_675_), .Y(_679_) );
	NOR2X1 NOR2X1_1145 ( .A(_672_), .B(_679_), .Y(_680_) );
	NOR3X1 NOR3X1_815 ( .A(_568_), .B(_588_), .C(_552_), .Y(_681_) );
	NOR3X1 NOR3X1_816 ( .A(_568_), .B(_588_), .C(_558_), .Y(_682_) );
	AOI22X1 AOI22X1_1527 ( .A(_681_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__0_), .D(_682_), .Y(_683_) );
	NOR3X1 NOR3X1_817 ( .A(_568_), .B(_582_), .C(_560_), .Y(_684_) );
	NOR3X1 NOR3X1_818 ( .A(_543_), .B(_553_), .C(_558_), .Y(_685_) );
	AOI22X1 AOI22X1_1528 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__0_), .B(_684_), .C(_685_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__0_), .Y(_686_) );
	NAND2X1 NAND2X1_2020 ( .A(_683_), .B(_686_), .Y(_687_) );
	NOR3X1 NOR3X1_819 ( .A(_582_), .B(_588_), .C(_568_), .Y(_688_) );
	NOR3X1 NOR3X1_820 ( .A(_558_), .B(_553_), .C(_572_), .Y(_689_) );
	AOI22X1 AOI22X1_1529 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__0_), .B(_688_), .C(_689_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__0_), .Y(_690_) );
	NOR3X1 NOR3X1_821 ( .A(_545_), .B(_553_), .C(_572_), .Y(_691_) );
	NOR3X1 NOR3X1_822 ( .A(_545_), .B(_588_), .C(_572_), .Y(_692_) );
	AOI22X1 AOI22X1_1530 ( .A(_691_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__0_), .D(_692_), .Y(_693_) );
	NAND2X1 NAND2X1_2021 ( .A(_693_), .B(_690_), .Y(_694_) );
	NOR2X1 NOR2X1_1146 ( .A(_687_), .B(_694_), .Y(_695_) );
	NAND2X1 NAND2X1_2022 ( .A(_695_), .B(_680_), .Y(_696_) );
	NOR3X1 NOR3X1_823 ( .A(_543_), .B(_582_), .C(_560_), .Y(_697_) );
	NOR3X1 NOR3X1_824 ( .A(_553_), .B(_562_), .C(_558_), .Y(_698_) );
	AOI22X1 AOI22X1_1531 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__0_), .B(_698_), .C(_697_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__0_), .Y(_699_) );
	NOR3X1 NOR3X1_825 ( .A(_547_), .B(_545_), .C(_572_), .Y(_700_) );
	NOR3X1 NOR3X1_826 ( .A(_558_), .B(_588_), .C(_572_), .Y(_701_) );
	AOI22X1 AOI22X1_1532 ( .A(_700_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__0_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__0_), .D(_701_), .Y(_702_) );
	NAND2X1 NAND2X1_2023 ( .A(_699_), .B(_702_), .Y(_703_) );
	NOR3X1 NOR3X1_827 ( .A(_543_), .B(_552_), .C(_560_), .Y(_704_) );
	NAND2X1 NAND2X1_2024 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__0_), .B(_704_), .Y(_705_) );
	NOR3X1 NOR3X1_828 ( .A(_562_), .B(_582_), .C(_547_), .Y(_706_) );
	NAND2X1 NAND2X1_2025 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__0_), .B(_706_), .Y(_707_) );
	NOR3X1 NOR3X1_829 ( .A(_545_), .B(_588_), .C(_568_), .Y(_708_) );
	NOR3X1 NOR3X1_830 ( .A(_545_), .B(_562_), .C(_560_), .Y(_709_) );
	AOI22X1 AOI22X1_1533 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__0_), .B(_708_), .C(_709_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__0_), .Y(_710_) );
	NAND3X1 NAND3X1_538 ( .A(_705_), .B(_707_), .C(_710_), .Y(_711_) );
	NOR2X1 NOR2X1_1147 ( .A(_711_), .B(_703_), .Y(_712_) );
	NOR3X1 NOR3X1_831 ( .A(_545_), .B(_568_), .C(_560_), .Y(_713_) );
	NOR3X1 NOR3X1_832 ( .A(_547_), .B(_562_), .C(_552_), .Y(_714_) );
	AOI22X1 AOI22X1_1534 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__0_), .B(_713_), .C(_714_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__0_), .Y(_715_) );
	NOR3X1 NOR3X1_833 ( .A(_547_), .B(_562_), .C(_558_), .Y(_716_) );
	NAND2X1 NAND2X1_2026 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__0_), .B(_716_), .Y(_717_) );
	NOR3X1 NOR3X1_834 ( .A(_552_), .B(_553_), .C(_572_), .Y(_718_) );
	NAND2X1 NAND2X1_2027 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__0_), .B(_718_), .Y(_719_) );
	NAND3X1 NAND3X1_539 ( .A(_717_), .B(_719_), .C(_715_), .Y(_720_) );
	NOR3X1 NOR3X1_835 ( .A(_552_), .B(_568_), .C(_560_), .Y(_721_) );
	NOR3X1 NOR3X1_836 ( .A(_562_), .B(_588_), .C(_545_), .Y(_722_) );
	AOI22X1 AOI22X1_1535 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__0_), .B(_722_), .C(_721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__0_), .Y(_723_) );
	NOR3X1 NOR3X1_837 ( .A(_558_), .B(_568_), .C(_560_), .Y(_724_) );
	NOR3X1 NOR3X1_838 ( .A(_562_), .B(_582_), .C(_553_), .Y(_725_) );
	AOI22X1 AOI22X1_1536 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__0_), .B(_725_), .C(_724_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__0_), .Y(_726_) );
	NAND2X1 NAND2X1_2028 ( .A(_723_), .B(_726_), .Y(_727_) );
	NOR2X1 NOR2X1_1148 ( .A(_727_), .B(_720_), .Y(_728_) );
	NAND2X1 NAND2X1_2029 ( .A(_712_), .B(_728_), .Y(_729_) );
	NOR3X1 NOR3X1_839 ( .A(_696_), .B(_665_), .C(_729_), .Y(_730_) );
	INVX1 INVX1_1240 ( .A(wSelec[13]), .Y(_731_) );
	NAND2X1 NAND2X1_2030 ( .A(wSelec[12]), .B(_731_), .Y(_732_) );
	INVX1 INVX1_1241 ( .A(wSelec[15]), .Y(_733_) );
	NAND2X1 NAND2X1_2031 ( .A(wSelec[14]), .B(_733_), .Y(_734_) );
	NOR2X1 NOR2X1_1149 ( .A(_732_), .B(_734_), .Y(_735_) );
	NOR2X1 NOR2X1_1150 ( .A(wSelec[13]), .B(wSelec[12]), .Y(_736_) );
	INVX1 INVX1_1242 ( .A(_736_), .Y(_737_) );
	NOR2X1 NOR2X1_1151 ( .A(_734_), .B(_737_), .Y(_738_) );
	AOI22X1 AOI22X1_1537 ( .A(wData[20]), .B(_735_), .C(_738_), .D(wData[16]), .Y(_739_) );
	INVX1 INVX1_1243 ( .A(wSelec[12]), .Y(_740_) );
	NAND2X1 NAND2X1_2032 ( .A(wSelec[13]), .B(_740_), .Y(_741_) );
	NOR2X1 NOR2X1_1152 ( .A(_741_), .B(_734_), .Y(_742_) );
	NAND2X1 NAND2X1_2033 ( .A(wData[24]), .B(_742_), .Y(_743_) );
	INVX1 INVX1_1244 ( .A(wSelec[14]), .Y(_744_) );
	NAND2X1 NAND2X1_2034 ( .A(_744_), .B(_733_), .Y(_745_) );
	NOR2X1 NOR2X1_1153 ( .A(_732_), .B(_745_), .Y(_746_) );
	NAND2X1 NAND2X1_2035 ( .A(wSelec[13]), .B(wSelec[12]), .Y(_747_) );
	NOR2X1 NOR2X1_1154 ( .A(_747_), .B(_734_), .Y(_748_) );
	AOI22X1 AOI22X1_1538 ( .A(_748_), .B(wData[28]), .C(wData[4]), .D(_746_), .Y(_749_) );
	NAND3X1 NAND3X1_540 ( .A(_743_), .B(_749_), .C(_739_), .Y(_750_) );
	NAND2X1 NAND2X1_2036 ( .A(wSelec[15]), .B(_744_), .Y(_751_) );
	NOR2X1 NOR2X1_1155 ( .A(_751_), .B(_737_), .Y(_752_) );
	NAND2X1 NAND2X1_2037 ( .A(wData[32]), .B(_752_), .Y(_753_) );
	NAND2X1 NAND2X1_2038 ( .A(wSelec[14]), .B(wSelec[15]), .Y(_754_) );
	NOR2X1 NOR2X1_1156 ( .A(_754_), .B(_741_), .Y(_755_) );
	NOR2X1 NOR2X1_1157 ( .A(_754_), .B(_732_), .Y(_756_) );
	AOI22X1 AOI22X1_1539 ( .A(_755_), .B(wData[56]), .C(wData[52]), .D(_756_), .Y(_757_) );
	NOR2X1 NOR2X1_1158 ( .A(_747_), .B(_754_), .Y(_758_) );
	NOR2X1 NOR2X1_1159 ( .A(_747_), .B(_751_), .Y(_759_) );
	AOI22X1 AOI22X1_1540 ( .A(wData[60]), .B(_758_), .C(_759_), .D(wData[44]), .Y(_760_) );
	NAND3X1 NAND3X1_541 ( .A(_753_), .B(_760_), .C(_757_), .Y(_761_) );
	NOR2X1 NOR2X1_1160 ( .A(_741_), .B(_751_), .Y(_762_) );
	NAND2X1 NAND2X1_2039 ( .A(wData[40]), .B(_762_), .Y(_763_) );
	NOR2X1 NOR2X1_1161 ( .A(_751_), .B(_732_), .Y(_764_) );
	NAND2X1 NAND2X1_2040 ( .A(wData[36]), .B(_764_), .Y(_765_) );
	NOR2X1 NOR2X1_1162 ( .A(_745_), .B(_737_), .Y(_766_) );
	NAND2X1 NAND2X1_2041 ( .A(wData[0]), .B(_766_), .Y(_767_) );
	NAND3X1 NAND3X1_542 ( .A(_763_), .B(_765_), .C(_767_), .Y(_768_) );
	INVX1 INVX1_1245 ( .A(wData[48]), .Y(_769_) );
	NOR2X1 NOR2X1_1163 ( .A(_744_), .B(_733_), .Y(_770_) );
	NAND2X1 NAND2X1_2042 ( .A(_736_), .B(_770_), .Y(_771_) );
	NOR2X1 NOR2X1_1164 ( .A(_741_), .B(_745_), .Y(_772_) );
	NOR2X1 NOR2X1_1165 ( .A(_747_), .B(_745_), .Y(_773_) );
	AOI22X1 AOI22X1_1541 ( .A(_772_), .B(wData[8]), .C(wData[12]), .D(_773_), .Y(_774_) );
	OAI21X1 OAI21X1_343 ( .A(_769_), .B(_771_), .C(_774_), .Y(_775_) );
	OR2X2 OR2X2_112 ( .A(_775_), .B(_768_), .Y(_776_) );
	NOR3X1 NOR3X1_840 ( .A(_750_), .B(_761_), .C(_776_), .Y(_777_) );
	AND2X2 AND2X2_214 ( .A(_777_), .B(_541_), .Y(_778_) );
	AOI21X1 AOI21X1_232 ( .A(_632_), .B(_730_), .C(_778_), .Y(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_0_) );
	INVX1 INVX1_1246 ( .A(_649_), .Y(_779_) );
	AOI21X1 AOI21X1_233 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__1_), .B(_779_), .C(_541_), .Y(_780_) );
	AOI22X1 AOI22X1_1542 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__1_), .B(_549_), .C(_565_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__1_), .Y(_781_) );
	AOI22X1 AOI22X1_1543 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__1_), .B(_569_), .C(_575_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__1_), .Y(_782_) );
	NAND3X1 NAND3X1_543 ( .A(_780_), .B(_781_), .C(_782_), .Y(_783_) );
	INVX1 INVX1_1247 ( .A(_609_), .Y(_784_) );
	AOI22X1 AOI22X1_1544 ( .A(_634_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__1_), .D(_784_), .Y(_785_) );
	AOI22X1 AOI22X1_1545 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__1_), .B(_708_), .C(_587_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__1_), .Y(_786_) );
	INVX1 INVX1_1248 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__1_), .Y(_787_) );
	INVX1 INVX1_1249 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__1_), .Y(_788_) );
	OAI22X1 OAI22X1_264 ( .A(_787_), .B(_596_), .C(_594_), .D(_788_), .Y(_789_) );
	INVX1 INVX1_1250 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__1_), .Y(_790_) );
	NAND2X1 NAND2X1_2043 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__1_), .B(_697_), .Y(_791_) );
	OAI21X1 OAI21X1_344 ( .A(_790_), .B(_602_), .C(_791_), .Y(_792_) );
	NOR2X1 NOR2X1_1166 ( .A(_789_), .B(_792_), .Y(_793_) );
	NAND3X1 NAND3X1_544 ( .A(_785_), .B(_786_), .C(_793_), .Y(_794_) );
	INVX1 INVX1_1251 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__1_), .Y(_795_) );
	NAND2X1 NAND2X1_2044 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__1_), .B(_581_), .Y(_796_) );
	OAI21X1 OAI21X1_345 ( .A(_795_), .B(_611_), .C(_796_), .Y(_797_) );
	INVX1 INVX1_1252 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__1_), .Y(_798_) );
	INVX1 INVX1_1253 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__1_), .Y(_799_) );
	OAI22X1 OAI22X1_265 ( .A(_798_), .B(_617_), .C(_615_), .D(_799_), .Y(_800_) );
	NOR2X1 NOR2X1_1167 ( .A(_800_), .B(_797_), .Y(_801_) );
	AOI22X1 AOI22X1_1546 ( .A(_701_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__1_), .D(_674_), .Y(_802_) );
	AND2X2 AND2X2_215 ( .A(_548_), .B(_563_), .Y(_803_) );
	AOI22X1 AOI22X1_1547 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__1_), .B(_673_), .C(_803_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__1_), .Y(_804_) );
	NAND3X1 NAND3X1_545 ( .A(_802_), .B(_804_), .C(_801_), .Y(_805_) );
	NOR3X1 NOR3X1_841 ( .A(_805_), .B(_783_), .C(_794_), .Y(_806_) );
	INVX1 INVX1_1254 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__1_), .Y(_807_) );
	NAND2X1 NAND2X1_2045 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__1_), .B(_636_), .Y(_808_) );
	OAI21X1 OAI21X1_346 ( .A(_638_), .B(_807_), .C(_808_), .Y(_809_) );
	AOI21X1 AOI21X1_234 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__1_), .B(_685_), .C(_809_), .Y(_810_) );
	INVX1 INVX1_1255 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__1_), .Y(_811_) );
	INVX1 INVX1_1256 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__1_), .Y(_812_) );
	OAI22X1 OAI22X1_266 ( .A(_812_), .B(_644_), .C(_645_), .D(_811_), .Y(_813_) );
	INVX1 INVX1_1257 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__1_), .Y(_814_) );
	NAND2X1 NAND2X1_2046 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__1_), .B(_654_), .Y(_815_) );
	OAI21X1 OAI21X1_347 ( .A(_555_), .B(_814_), .C(_815_), .Y(_816_) );
	NOR2X1 NOR2X1_1168 ( .A(_816_), .B(_813_), .Y(_817_) );
	INVX1 INVX1_1258 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__1_), .Y(_818_) );
	INVX1 INVX1_1259 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__1_), .Y(_819_) );
	OAI22X1 OAI22X1_267 ( .A(_650_), .B(_819_), .C(_656_), .D(_818_), .Y(_820_) );
	INVX1 INVX1_1260 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__1_), .Y(_821_) );
	NOR2X1 NOR2X1_1169 ( .A(_821_), .B(_661_), .Y(_822_) );
	INVX1 INVX1_1261 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__1_), .Y(_823_) );
	NOR2X1 NOR2X1_1170 ( .A(_823_), .B(_662_), .Y(_824_) );
	NOR3X1 NOR3X1_842 ( .A(_822_), .B(_820_), .C(_824_), .Y(_825_) );
	NAND3X1 NAND3X1_546 ( .A(_817_), .B(_810_), .C(_825_), .Y(_826_) );
	AOI22X1 AOI22X1_1548 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__1_), .B(_666_), .C(_667_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__1_), .Y(_827_) );
	AOI22X1 AOI22X1_1549 ( .A(_669_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__1_), .D(_670_), .Y(_828_) );
	NAND2X1 NAND2X1_2047 ( .A(_827_), .B(_828_), .Y(_829_) );
	AOI22X1 AOI22X1_1550 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__1_), .B(_677_), .C(_676_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__1_), .Y(_830_) );
	AOI22X1 AOI22X1_1551 ( .A(_620_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__1_), .D(_627_), .Y(_831_) );
	NAND2X1 NAND2X1_2048 ( .A(_830_), .B(_831_), .Y(_832_) );
	NOR2X1 NOR2X1_1171 ( .A(_829_), .B(_832_), .Y(_833_) );
	AOI22X1 AOI22X1_1552 ( .A(_681_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__1_), .D(_682_), .Y(_834_) );
	AOI22X1 AOI22X1_1553 ( .A(_583_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__1_), .D(_684_), .Y(_835_) );
	NAND2X1 NAND2X1_2049 ( .A(_834_), .B(_835_), .Y(_836_) );
	AOI22X1 AOI22X1_1554 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__1_), .B(_688_), .C(_689_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__1_), .Y(_837_) );
	AOI22X1 AOI22X1_1555 ( .A(_691_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__1_), .D(_692_), .Y(_838_) );
	NAND2X1 NAND2X1_2050 ( .A(_838_), .B(_837_), .Y(_839_) );
	NOR2X1 NOR2X1_1172 ( .A(_836_), .B(_839_), .Y(_840_) );
	NAND2X1 NAND2X1_2051 ( .A(_840_), .B(_833_), .Y(_841_) );
	AOI22X1 AOI22X1_1556 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__1_), .B(_698_), .C(_599_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__1_), .Y(_842_) );
	AOI22X1 AOI22X1_1557 ( .A(_622_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__1_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__1_), .D(_700_), .Y(_843_) );
	NAND2X1 NAND2X1_2052 ( .A(_842_), .B(_843_), .Y(_844_) );
	AOI22X1 AOI22X1_1558 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__1_), .B(_589_), .C(_709_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__1_), .Y(_845_) );
	NAND2X1 NAND2X1_2053 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__1_), .B(_704_), .Y(_846_) );
	NAND2X1 NAND2X1_2054 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__1_), .B(_706_), .Y(_847_) );
	NAND3X1 NAND3X1_547 ( .A(_846_), .B(_847_), .C(_845_), .Y(_848_) );
	NOR2X1 NOR2X1_1173 ( .A(_848_), .B(_844_), .Y(_849_) );
	AOI22X1 AOI22X1_1559 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__1_), .B(_713_), .C(_714_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__1_), .Y(_850_) );
	NAND2X1 NAND2X1_2055 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__1_), .B(_716_), .Y(_851_) );
	NAND2X1 NAND2X1_2056 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__1_), .B(_718_), .Y(_852_) );
	NAND3X1 NAND3X1_548 ( .A(_851_), .B(_852_), .C(_850_), .Y(_853_) );
	AOI22X1 AOI22X1_1560 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__1_), .B(_722_), .C(_721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__1_), .Y(_854_) );
	AOI22X1 AOI22X1_1561 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__1_), .B(_725_), .C(_724_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__1_), .Y(_855_) );
	NAND2X1 NAND2X1_2057 ( .A(_854_), .B(_855_), .Y(_856_) );
	NOR2X1 NOR2X1_1174 ( .A(_856_), .B(_853_), .Y(_857_) );
	NAND2X1 NAND2X1_2058 ( .A(_849_), .B(_857_), .Y(_858_) );
	NOR3X1 NOR3X1_843 ( .A(_841_), .B(_826_), .C(_858_), .Y(_859_) );
	AOI21X1 AOI21X1_235 ( .A(wData[21]), .B(_735_), .C(_540_), .Y(_860_) );
	AOI22X1 AOI22X1_1562 ( .A(_738_), .B(wData[17]), .C(wData[1]), .D(_766_), .Y(_861_) );
	AOI22X1 AOI22X1_1563 ( .A(_759_), .B(wData[45]), .C(wData[25]), .D(_742_), .Y(_862_) );
	NAND3X1 NAND3X1_549 ( .A(_860_), .B(_862_), .C(_861_), .Y(_863_) );
	NAND3X1 NAND3X1_550 ( .A(wData[49]), .B(_736_), .C(_770_), .Y(_864_) );
	AOI22X1 AOI22X1_1564 ( .A(wData[61]), .B(_758_), .C(_746_), .D(wData[5]), .Y(_865_) );
	AND2X2 AND2X2_216 ( .A(_865_), .B(_864_), .Y(_866_) );
	AOI22X1 AOI22X1_1565 ( .A(_755_), .B(wData[57]), .C(wData[41]), .D(_762_), .Y(_867_) );
	AOI22X1 AOI22X1_1566 ( .A(wData[53]), .B(_756_), .C(_752_), .D(wData[33]), .Y(_868_) );
	AND2X2 AND2X2_217 ( .A(_868_), .B(_867_), .Y(_869_) );
	AOI22X1 AOI22X1_1567 ( .A(_772_), .B(wData[9]), .C(wData[13]), .D(_773_), .Y(_870_) );
	AOI22X1 AOI22X1_1568 ( .A(_748_), .B(wData[29]), .C(wData[37]), .D(_764_), .Y(_871_) );
	AND2X2 AND2X2_218 ( .A(_870_), .B(_871_), .Y(_872_) );
	NAND3X1 NAND3X1_551 ( .A(_866_), .B(_872_), .C(_869_), .Y(_873_) );
	NOR2X1 NOR2X1_1175 ( .A(_863_), .B(_873_), .Y(_874_) );
	AOI21X1 AOI21X1_236 ( .A(_806_), .B(_859_), .C(_874_), .Y(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_1_) );
	AOI21X1 AOI21X1_237 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__2_), .B(_779_), .C(_541_), .Y(_875_) );
	INVX1 INVX1_1262 ( .A(_638_), .Y(_876_) );
	AOI22X1 AOI22X1_1569 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__2_), .B(_549_), .C(_876_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__2_), .Y(_877_) );
	INVX1 INVX1_1263 ( .A(_650_), .Y(_878_) );
	AOI22X1 AOI22X1_1570 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_18__2_), .B(_685_), .C(_878_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__2_), .Y(_879_) );
	NAND3X1 NAND3X1_552 ( .A(_879_), .B(_875_), .C(_877_), .Y(_880_) );
	AOI22X1 AOI22X1_1571 ( .A(_634_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__2_), .D(_784_), .Y(_881_) );
	AOI22X1 AOI22X1_1572 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__2_), .B(_583_), .C(_556_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__2_), .Y(_882_) );
	INVX1 INVX1_1264 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__2_), .Y(_883_) );
	NAND2X1 NAND2X1_2059 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_40__2_), .B(_673_), .Y(_884_) );
	OAI21X1 OAI21X1_348 ( .A(_883_), .B(_645_), .C(_884_), .Y(_885_) );
	INVX1 INVX1_1265 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__2_), .Y(_886_) );
	NAND2X1 NAND2X1_2060 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_26__2_), .B(_599_), .Y(_887_) );
	OAI21X1 OAI21X1_349 ( .A(_886_), .B(_602_), .C(_887_), .Y(_888_) );
	NOR2X1 NOR2X1_1176 ( .A(_885_), .B(_888_), .Y(_889_) );
	NAND3X1 NAND3X1_553 ( .A(_881_), .B(_882_), .C(_889_), .Y(_890_) );
	INVX1 INVX1_1266 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__2_), .Y(_891_) );
	NAND2X1 NAND2X1_2061 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__2_), .B(_581_), .Y(_892_) );
	OAI21X1 OAI21X1_350 ( .A(_891_), .B(_611_), .C(_892_), .Y(_893_) );
	INVX1 INVX1_1267 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__2_), .Y(_894_) );
	INVX1 INVX1_1268 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__2_), .Y(_895_) );
	OAI22X1 OAI22X1_268 ( .A(_894_), .B(_617_), .C(_615_), .D(_895_), .Y(_896_) );
	NOR2X1 NOR2X1_1177 ( .A(_896_), .B(_893_), .Y(_897_) );
	AOI22X1 AOI22X1_1573 ( .A(_701_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_46__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_41__2_), .D(_674_), .Y(_898_) );
	AND2X2 AND2X2_219 ( .A(_573_), .B(_595_), .Y(_899_) );
	AOI22X1 AOI22X1_1574 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__2_), .B(_899_), .C(_803_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_52__2_), .Y(_900_) );
	NAND3X1 NAND3X1_554 ( .A(_898_), .B(_900_), .C(_897_), .Y(_901_) );
	NOR3X1 NOR3X1_844 ( .A(_901_), .B(_880_), .C(_890_), .Y(_902_) );
	INVX1 INVX1_1269 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_1__2_), .Y(_903_) );
	NOR3X1 NOR3X1_845 ( .A(_903_), .B(_568_), .C(_567_), .Y(_904_) );
	AND2X2 AND2X2_220 ( .A(_589_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_63__2_), .Y(_905_) );
	AND2X2 AND2X2_221 ( .A(_709_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_56__2_), .Y(_906_) );
	NOR3X1 NOR3X1_846 ( .A(_906_), .B(_905_), .C(_904_), .Y(_907_) );
	INVX1 INVX1_1270 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_57__2_), .Y(_908_) );
	INVX1 INVX1_1271 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_28__2_), .Y(_909_) );
	OAI22X1 OAI22X1_269 ( .A(_909_), .B(_644_), .C(_594_), .D(_908_), .Y(_910_) );
	INVX1 INVX1_1272 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_58__2_), .Y(_911_) );
	INVX1 INVX1_1273 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_2__2_), .Y(_912_) );
	NAND2X1 NAND2X1_2062 ( .A(_585_), .B(_586_), .Y(_913_) );
	OAI22X1 OAI22X1_270 ( .A(_913_), .B(_912_), .C(_911_), .D(_564_), .Y(_914_) );
	NOR2X1 NOR2X1_1178 ( .A(_910_), .B(_914_), .Y(_915_) );
	INVX1 INVX1_1274 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_37__2_), .Y(_916_) );
	NOR3X1 NOR3X1_847 ( .A(_545_), .B(_562_), .C(_553_), .Y(_917_) );
	NAND2X1 NAND2X1_2063 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_48__2_), .B(_917_), .Y(_918_) );
	OAI21X1 OAI21X1_351 ( .A(_574_), .B(_916_), .C(_918_), .Y(_919_) );
	INVX1 INVX1_1275 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_49__2_), .Y(_920_) );
	INVX1 INVX1_1276 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_30__2_), .Y(_921_) );
	OAI22X1 OAI22X1_271 ( .A(_661_), .B(_921_), .C(_920_), .D(_662_), .Y(_922_) );
	NOR2X1 NOR2X1_1179 ( .A(_919_), .B(_922_), .Y(_923_) );
	NAND3X1 NAND3X1_555 ( .A(_907_), .B(_923_), .C(_915_), .Y(_924_) );
	AOI22X1 AOI22X1_1575 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_0__2_), .B(_666_), .C(_667_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_61__2_), .Y(_925_) );
	AOI22X1 AOI22X1_1576 ( .A(_669_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_62__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_59__2_), .D(_670_), .Y(_926_) );
	NAND2X1 NAND2X1_2064 ( .A(_925_), .B(_926_), .Y(_927_) );
	AOI22X1 AOI22X1_1577 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_31__2_), .B(_677_), .C(_676_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_29__2_), .Y(_928_) );
	AOI22X1 AOI22X1_1578 ( .A(_620_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_45__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_42__2_), .D(_627_), .Y(_929_) );
	NAND2X1 NAND2X1_2065 ( .A(_928_), .B(_929_), .Y(_930_) );
	NOR2X1 NOR2X1_1180 ( .A(_927_), .B(_930_), .Y(_931_) );
	AOI22X1 AOI22X1_1579 ( .A(_681_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_13__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_14__2_), .D(_682_), .Y(_932_) );
	AOI22X1 AOI22X1_1580 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_12__2_), .B(_708_), .C(_684_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_11__2_), .Y(_933_) );
	NAND2X1 NAND2X1_2066 ( .A(_933_), .B(_932_), .Y(_934_) );
	AOI22X1 AOI22X1_1581 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_15__2_), .B(_688_), .C(_689_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_34__2_), .Y(_935_) );
	AOI22X1 AOI22X1_1582 ( .A(_691_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_32__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_44__2_), .D(_692_), .Y(_936_) );
	NAND2X1 NAND2X1_2067 ( .A(_936_), .B(_935_), .Y(_937_) );
	NOR2X1 NOR2X1_1181 ( .A(_934_), .B(_937_), .Y(_938_) );
	NAND2X1 NAND2X1_2068 ( .A(_938_), .B(_931_), .Y(_939_) );
	AOI22X1 AOI22X1_1583 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_50__2_), .B(_698_), .C(_697_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__2_), .Y(_940_) );
	AOI22X1 AOI22X1_1584 ( .A(_622_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_43__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_36__2_), .D(_700_), .Y(_941_) );
	NAND2X1 NAND2X1_2069 ( .A(_940_), .B(_941_), .Y(_942_) );
	AOI22X1 AOI22X1_1585 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_55__2_), .B(_706_), .C(_704_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_25__2_), .Y(_943_) );
	AOI22X1 AOI22X1_1586 ( .A(_636_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_4__2_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__2_), .D(_654_), .Y(_944_) );
	NAND2X1 NAND2X1_2070 ( .A(_944_), .B(_943_), .Y(_945_) );
	NOR2X1 NOR2X1_1182 ( .A(_945_), .B(_942_), .Y(_946_) );
	AOI22X1 AOI22X1_1587 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_8__2_), .B(_713_), .C(_714_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_53__2_), .Y(_947_) );
	NAND2X1 NAND2X1_2071 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_54__2_), .B(_716_), .Y(_948_) );
	NAND2X1 NAND2X1_2072 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_33__2_), .B(_718_), .Y(_949_) );
	NAND3X1 NAND3X1_556 ( .A(_948_), .B(_949_), .C(_947_), .Y(_950_) );
	AOI22X1 AOI22X1_1588 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_60__2_), .B(_722_), .C(_721_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_9__2_), .Y(_951_) );
	AOI22X1 AOI22X1_1589 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_51__2_), .B(_725_), .C(_724_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_10__2_), .Y(_952_) );
	NAND2X1 NAND2X1_2073 ( .A(_951_), .B(_952_), .Y(_953_) );
	NOR2X1 NOR2X1_1183 ( .A(_953_), .B(_950_), .Y(_954_) );
	NAND2X1 NAND2X1_2074 ( .A(_946_), .B(_954_), .Y(_955_) );
	NOR3X1 NOR3X1_848 ( .A(_939_), .B(_924_), .C(_955_), .Y(_956_) );
	AOI22X1 AOI22X1_1590 ( .A(_762_), .B(wData[42]), .C(wData[38]), .D(_764_), .Y(_957_) );
	AOI22X1 AOI22X1_1591 ( .A(_759_), .B(wData[46]), .C(_766_), .D(wData[2]), .Y(_958_) );
	NAND2X1 NAND2X1_2075 ( .A(_957_), .B(_958_), .Y(_959_) );
	AOI21X1 AOI21X1_238 ( .A(wData[34]), .B(_752_), .C(_959_), .Y(_960_) );
	INVX1 INVX1_1277 ( .A(wData[50]), .Y(_961_) );
	AOI22X1 AOI22X1_1592 ( .A(_772_), .B(wData[10]), .C(wData[14]), .D(_773_), .Y(_962_) );
	OAI21X1 OAI21X1_352 ( .A(_961_), .B(_771_), .C(_962_), .Y(_963_) );
	AOI22X1 AOI22X1_1593 ( .A(_735_), .B(wData[22]), .C(wData[18]), .D(_738_), .Y(_964_) );
	NAND2X1 NAND2X1_2076 ( .A(wData[26]), .B(_742_), .Y(_965_) );
	AOI22X1 AOI22X1_1594 ( .A(_748_), .B(wData[30]), .C(wData[6]), .D(_746_), .Y(_966_) );
	NAND3X1 NAND3X1_557 ( .A(_965_), .B(_966_), .C(_964_), .Y(_967_) );
	NOR2X1 NOR2X1_1184 ( .A(_963_), .B(_967_), .Y(_968_) );
	NAND2X1 NAND2X1_2077 ( .A(wData[58]), .B(_755_), .Y(_969_) );
	NAND2X1 NAND2X1_2078 ( .A(wData[54]), .B(_756_), .Y(_970_) );
	NAND2X1 NAND2X1_2079 ( .A(_969_), .B(_970_), .Y(_971_) );
	AOI21X1 AOI21X1_239 ( .A(wData[62]), .B(_758_), .C(_971_), .Y(_972_) );
	NAND3X1 NAND3X1_558 ( .A(_960_), .B(_972_), .C(_968_), .Y(_973_) );
	NOR2X1 NOR2X1_1185 ( .A(_540_), .B(_973_), .Y(_974_) );
	AOI21X1 AOI21X1_240 ( .A(_902_), .B(_956_), .C(_974_), .Y(input_selector_block_input_selector_i_0__input_selector_j_1__input_selector_r_2_) );
	AOI21X1 AOI21X1_241 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_22__3_), .B(_784_), .C(_541_), .Y(_975_) );
	AOI22X1 AOI22X1_1595 ( .A(_556_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_17__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_6__3_), .D(_876_), .Y(_976_) );
	AOI22X1 AOI22X1_1596 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_3__3_), .B(_878_), .C(_634_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_23__3_), .Y(_977_) );
	NAND3X1 NAND3X1_559 ( .A(_977_), .B(_975_), .C(_976_), .Y(_978_) );
	AOI22X1 AOI22X1_1597 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_19__3_), .B(_583_), .C(_581_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_16__3_), .Y(_979_) );
	AOI22X1 AOI22X1_1598 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_7__3_), .B(_654_), .C(_779_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_21__3_), .Y(_980_) );
	INVX1 INVX1_1278 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_47__3_), .Y(_981_) );
	INVX1 INVX1_1279 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_5__3_), .Y(_982_) );
	OAI22X1 OAI22X1_272 ( .A(_981_), .B(_596_), .C(_645_), .D(_982_), .Y(_983_) );
	INVX1 INVX1_1280 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_39__3_), .Y(_984_) );
	NAND2X1 NAND2X1_2080 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_27__3_), .B(_697_), .Y(_985_) );
	OAI21X1 OAI21X1_353 ( .A(_984_), .B(_602_), .C(_985_), .Y(_986_) );
	NOR2X1 NOR2X1_1186 ( .A(_983_), .B(_986_), .Y(_987_) );
	NAND3X1 NAND3X1_560 ( .A(_979_), .B(_980_), .C(_987_), .Y(_988_) );
	AND2X2 AND2X2_222 ( .A(_610_), .B(_544_), .Y(_989_) );
	AOI22X1 AOI22X1_1599 ( .A(_549_), .B(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_20__3_), .C(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_24__3_), .D(_989_), .Y(_990_) );
	AND2X2 AND2X2_223 ( .A(_608_), .B(_573_), .Y(_991_) );
	AND2X2 AND2X2_224 ( .A(_616_), .B(_573_), .Y(_992_) );
	AOI22X1 AOI22X1_1600 ( .A(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_35__3_), .B(_992_), .C(_991_), .D(input_selector_block_input_selector_i_0__input_selector_j_0__input_selector_chunksRegs_38__3_), .Y(_993_) );
endmodule
